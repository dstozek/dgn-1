��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-?H)t� �hz2��ƿ� �lJE�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hp���Ť�Mn��X)r����#�L������5N�1 T�V	�tL��	�{�Κ$M�C7y���v6޿���kq����Eֿ�o0��ܧe���5�/���ׇӭ��!�`�(i3[�"5�QJǊö��_��i@�{ۧe[ғr�,�Ōt�}Uٱ�g����.E�^~_|�����{j�G:� ��'��iI+w,A��4�M\���Z ��a�O>*���
��#kz��GN�P�0v���uP!ߌ���^����Wړ��]b�=#;6�#t����nB3�+{Cz��3�<A��d�]��<��&�gG��Hc�e$���=�(v
���O>E$I������T���Q���!i��ӯ�0���&�:�u0&����x2�Zy����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�jM�1}2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!����j.�n�Ax��PR@?�Q|33�����rqn���wѪ	/g�%�W��{�RX�>w�P���u0�������k�V�99^�)�S��uC|Q�����9�ih\���6�oX��s�At�Ӡ�-������u�=�xs�1����";1�(�����]a�{��ۊ�d�k�`�?��<�� ��o�}a�Còz�;^�ru��e��_$߼
�d�YiUbiX>�"��g��3�G��/8'��ި]M�}xf���T��Mߟy�����n��1��\�p��/L�M��Y�Ҁ����r��{��>ڑ/8'�odgƚ�| �����q��5k�^�78���N��ov�Op����	�Y8�>����;% ���W~�_Y�1�����q[��\�jf)�bdZ0o�v�v���O��q�M�4��{i�etWj%h�W�8������8ٓ�j!�`�(i3p]G��>���<�}��x~QTߨ�O3��\�'�y'��BS�z�5&n��ū��@�k�!�`�(i3!�`�(i3!�`�(i3}[x��8��`��Ć?6�!s}6,e �ǟ=EZئ;z&����+�E�r{����JDn ��a�K�.:gdW(o%�)���;t|������D"�~����p�4���='߰����`H��b/3j!�`�(i3!�`�(i3�F{/���!3~�(Z��GmO��%��}�.����M���5^s1@�&'iKb�آ[�~,ΗG\�ʢ�X�=1�����
�^��j"��Q�]f�p����=Qsz����Iv�.�GzEc.������������X�k=o���Fz�!�`�(i3!�`�(i3IB�]�!P���b6p!!v*!���&fB�@��X*,l��d���F6���ׇӭ��!�`�(i3!�`�(i3 lF�Z��f}�y�F�&��S߭;�(6��3{��|o	���=l"�,�>E��&�3�y�2��J�J�T�S1(_�'�&r�~,ptQ��k$Vʴ8X�S����TXP�e�g]�H��֟B��Ўek'`�j�13*�á)ˎ	��[�!%&oA�\ֆ�
'��(�<��
Aʎ^g!�`�(i3!�`�(i3!�`�(i3�|j��"C���ޝsn?V��-Q	�	:����lg\ ����EO�{��ϫ��u�o���q�Z��?��: 0[�T#�l�/Zw������{%hPb��͓T�)��z��z
��K�O�n���^���D�*�Z�J�v$��A�f�y'��BSƹ�#�y�w���	B$�@�A�w{6��(�N��K�O�n8�[ �n�
�CQYb!��uፁ�&�$`8�+DO�n�;4L&�y;U�2y��}���[N�)J��7)�c�0:S��}1yYZ��� ����@	�1i�myh�~�*�.i,����j�Ə���&,���9�tOHn����x���I8I�%-4o��Iu���'�#&��
 {�L<��-�|��e���RB����bb��Ə���&,��+���!XwOHn����x���I8I�%-4o��Iu���'�#&_�:q`��� �Z)}�6!ת���ېư���o���o��V�x�O`BpI�ҽb.j����kѶ���� ���X%��m�Z9a\������0;8�y�%$���r���{��6;)ܟaTo0BpI�ҽb.j����#�2�/D<�L�k��\|�M4��*��J�Y��в}��aC�2V�Vׇӭ��!�`�(i3!�`�(i3I����Ǻ'n;�>�rY
�����+O~%��짐~��.d����"���p|��X^䀸~�W߁�nrm؊(�[���~$�B2���m���-��
�8���?�*���\�Ə���&,Ƿ	DTjE,���6��q@�2��>�b!��u�Z1~�g]�u�+��
~J[����30�A�zc�RhoŜn!�`�(i3!�`�(i3!�`�(i3�M��n���<����lpU�:�ƅf��	��������6��q@�2��>�o����|�sg�2�:��~�^=��D�,<�V�QK�}�9���u����Fz�!�`�(i3!�`�(i3؝�4W���+DO�n��t!I����;R���fǥ�c⠵���طYRdZ0o�v�V#��ب'�����{��6;<� ֭m�_���ȃEE��$(��{�$�˽�Lk�`�?��<��t!I������h+�w��4܆��O�2C��OG;�['*�p!!v*!���O�{�
;����"����+H]�����˶���,/Pc��?@W��8�����b2�{������7��U�:�ƅf�H��������6�����+��w-���f*���׎o�|��Y�� �k��^��Xz�Ȗ��W�{N������~چ�sֱ"MT}���o�׎o�|��Y�� �k��^��Xz�(��¦�L\�kg�Ť����� E��5�O�U���.b!��u�w���v.���A�I�z�9w+�!J�0©	]�,�\DW.ɧ/H>y7�J�]f7\��1�T�g��������G2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcn��^��N�oߛN�N�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hF^����i�̨���qh�'aba�	���
��?��n;�|-�Z��2S ���k��m���$[΁�a�n��Vk��w/&g�-ΘBdN�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_c9��*��OT��]S��f����om2�����iҢ��V�x��%�a��i�9�J��$b6�]ʆ�In��t@���z������)����")�^�3��8r�Wk�ǻow��R�nI�GI$��ǂcY�~遅��'�:��'n�^0o��S��S�Ib���ό���.ӥóM�˄NQ��臿5"c'��ɿ��3P�d�8!��vp�P}��O���w2T��b�T��xd�Y�I�;\h!E��c�G�*ZkS0��nB�+������]��)`���"��y�LN��K��g����R�<�W�C%c�����<�W�C%����_Wr��;���EWr�L{1��ox ������ �i7�sp>{=J���.��W�}�"�,�>E����\�vūx`��:��g�0�u�L{1��oxr�O΅��C?�D�s�R�"0��<��	��������JF!՟Ր��M�aW��Σ�?��<��z�"�~��S�
/P��Ѷ����A5wr�4�Vgn`��p���n�O�V�N�s
l���u���NX@��^��>��}� ���O%��y�䃶&f�����SVc�5ߧE4��?"����a�m���q�l;1�]�I�rT�8#�>-��;��S������yq]C
R��T
�N�oߛN�N�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hF^����i�̨���qh�'aba�	���
��?��n;�|-�Z��2S ���k��m���$[΁�a�n��Vk��w/&g�-ΘBdN�FQx�0O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_c9��*��OT��]S��f����om2�n�h޶�\�Ji��'�o��Q$������aU��D�	a���(�E��!�`�(i3l0��F��j���^B_�(ba�7�X��)z�s�!�`�(i3%Ah�%4
>��XP��Ȱ�^�7^/�AJy���l�f�nϵ ���3�ҺIÙ=�H�}ʧ8Еb����������gE�,�Q�^�y�zL͊�q��_�0���ӨI��'���Z[A�E����F�'n�^0oL��pN�5����`K�x��R͖"�,�>E����\�vŻA�1�#`�͌4s+�ny���A�!3v!�`�(i3JHn��z� �&�^`(���%�a�N�+��#�!�`�(i3�b9���6,� k\\1�*_��hc�ʹ���`!�`�(i3l0��F��j���^B_�||�?�5���J��xi��͆'�X%Ah�%4
>��XP��ȵ�d��w����y{¦�$]\� ���3�ҺIÙ=�H�uoglR���c&;�p� ���S�Q�^�y�zL͊�q�� �-8���I��'�	�ų_��E����F�'n�^0o%|�J�0�5����`K��q��"�,�>E����\�v�Qq
˟6͌4s+�ny��9� W0�!�`�(i3JHn��z�k��%��6i��%�a�x�+Vv��2!�`�(i3�b9���
Ay�9�6>1�*_��h���Q��~��
c�[��ƣD��T�����NI�����m�2�Z,qC͌4s+�nycfl��6t�$X4P�JHn��z�S@�z�R3��%�a������?6�9������7s�9���o��S8��%�CF�I��r��Ȯ��ߊ��H�R�?�ɺdX�-�B�85���%�a������?6E�C�Έ��7s�9���o��S8��%�CF�I��r��Ȯ��ߊ��H�R�?�ɺdX��<�-���#�p������p:�2],˶�9�c	o'E!��s�Zu�EPD]�I���2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p���}������]�0�lK'���Xw��_
�u�m�\��q�Z˻r������U�r�}��}����ހmu�m����y^�k���%H�$N�oߛN�cL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!��D���X=��f��i��зq8�ЈxKʜ�#xI+r�� 0�D�A��t��D)��i�d��`m�¨3��%�$�������\O�a�|�6����&��DErwⳘ=�C. ��f?��s^�xct��_Tҥ!�V��NR0�����O�,�WNT�N D|�5N��VA}�v�a'����\�Z��'�Wa�L��ʻR0�˧���.�E����Fr<���\�g�-ΘBdcL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U��k�t���L53�����)-}�vPt�>xA�ꓩ�l;��!I/�������A��1��+�W��J�ݨg4$ _o����OI��@���:��F�b��@�zL͊�q��c�sYIJ8��OI��@�n���������Wq{�f��a��{oS�=wK��7�&d&(C�#�7#^�Vn�^ֻ����XP��Ȇ<�qp^S��j.Z��$�sӢ�]3�����c��(r$����G���'aOދK-\��$-��Ǡ٥L����e]�u�����!�M�T���ݏ��A�!�`�(i3���+�J�������"�,�>E��W��Ґ�YjZ�p��Z����r;��*!�`�(i3"�,�>E����\�v�!�`�(i3Sn<Z�)K|K�@�����!�+�!�`�(i3%Ah�%4
>��f���T,�;C@����%?!m�Az�F��O�4p���eq��VZ�0�s�b<�B�_���X�KM�����7������
�]qE�&���W����Q�^�y�����9�!�`�(i3���3�b���-the��戉Z�T!�`�(i37s�9���o��S8����J� �j��h@S�@�]_LO!�`�(i3JHn��z��x�f7﹏�1β��h����0���,�W�B�޹B$~s%��@�:�����xwƄ�{Ƨ\-TX�Rj�+s�!���r��*y�xDp��T�/i�M���"�,�>E����\�v�!�`�(i3y�Er�)=�ᏅN~z��9�{�G�K*V׹ږ��_��f���T,�;C@����P@zQX�76�$t8[��5��FX9�p�x^/8�D�n�ؒ1ECWI�R��R��=���b>���F9M؛��&�}�(�dW�,��(�a�肢�{l�f|�ό���.ӟ
�r��	G$��R�lD<��z��}�Q2�+�Yə~�yD݃��r��DB�����I�b}Ω:���V�(^��<��z��}�Q2�+�Y�7
�4�.�E����F�ҋX����|P�������A�=�8bH���L��B�;#5d���7Ê7�E�4'���Xw/���:;aR[�T�.�W���1�}�ױ��(@�E����F�ҋX����|P�������A�=�8bH���L��B��)�ޭ-�7Ê7�E�4'���Xw/���:;aR[�T�.�W���1��)$磨'jU-j�`�ҋX����|P�������A�=�8bH��Ę媌�+�<1(f}ظ{����$ <��HT� \r���㯄�����
L'���Xw��RN�-#�ьb2up,zk�g��[��v�$ƪ;���Q��/(A=�kX�*1�e38����2�9)�����m��T��J<�]qE�&�owђN�~R�wX�յ�8�,wO۳�yz�<��z��}�0z�cUL� ���Q�'e����u*w�A	'���k(�պ6<��z��}�0z�cUL� ���Q�'e����-��\4vߖ%��mz%���=a\�&'UR�q������3���R����o秾�!a�v�����w:ꮆ@IE�U��@�ڗe'a�v�����*� ���@IE�U��@�ڗe'����h+������E��@IE�U��@�ڗe'��;R����H���i�Ox�j�d�ƥ4�,�:�'t��t�W�lT[�HF x>H�|�Wǖg3ȓ8���/�A���0v7���V�x�O`�����
L'���Xw�j�7���rcJ]�0ݫ���Uh1�gؘC���t\>��fm��]2�y�Z鎬����)��e���Rf?����]2�y�Z鎬����)��e���= �J4��]2�y�Z鎬����L�`u�K�˱�Ui��Q�x��8�,wO��ٷ���TD��-�`��8�4�%��mz%���=a\�9�K�v`0���'=��"B��$I��w��,��xc�l��m
��5�(�����:x�V?W�)�ޭ-����
L'���Xw/���:;aR[�T�.�W���1���~������yf��?N/7G#+������z����A�b�*܋���ԓ�Dd�<�,E9|.���%�S��v���?�R����o秾�!rF)���X�3c/��!ő!XF3�@IE�U��@�ڗe'rF)���X�3c/��!�:GV��d@@IE�U��@�ڗe'rF)���X�3c/��!P;��	�@IE�U��@�ڗe'rF)���X�3c/��!4V(�x@IE�U��@�ڗe'rF)���X�3c/��!з���jf@IE�U��@�ڗe'rF)���X�3c/��!�f���l @IE�U��@�ڗe'rF)���X�3c/��!�Q��Y��@IE�U��@�ڗe'rF)���X�3c/��!��8�ۦ@IE�U��@�ڗe'rF)���X�3c/��!��A Ly�@IE�U��@�ڗe'rF)���X�3c/��!k�O�`c @IE�U��@�ڗe'rF)���X�3c/��!����4��8@IE�U��@�ڗe'rF)���X�3c/��!.�0�;l@IE�U��@�ڗe'rF)���X�3c/��!'��t#~t@IE�U��@�ڗe'rF)���X�3c/��!򊫖��@IE�U��@�ڗe'rF)���X�3c/��!��];p��@IE�U��@�ڗe'rF)���X�3c/��!���L���@IE�U��*�QN��� ]���f��v�鳔�Ċ��8���K(��z�j�;9�e��L53���Z<�~�q��]3�����c��(r�CRQ���E�+d�ίp��V�����Y����딼�\�v���T�©�#��l�َ2c�'z͌4s+�ny�X��{��ܛ�	�����^�%k IÙ=�Ho?Y���	3�Ð�9�X�e�B���<����ą~c�PƐt
����������\�v���T�©@���U@���:��F�����XuY*"�nw��F�dZ0o�v��CRQ���Eu<�.��	�L�t0{�A����8V�l0��F��j.��h��u>1�*_��h��Ӯw!)��&�t5C�,���m�b9������U.6����sd�Hc�.2��w�k#�J����͌4s+�ny\D}��^�y�����"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s�6F���y�8� �w� G�"�|� }�Ri.����l���r{����JDn ��aů�x� ���rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'��KD����w�Ve�U�ԝ5�͌4s+�ny7\�%Lţ}���u=|�z�)�]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s���A0�>�8� �w� G�"�|� }�Ri.����l���R�0�;"��9�{���|hY���rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'��QV&�f�w�Ve�U�ԝ5�͌4s+�ny�y��P�p�V��O"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��{_8�Y���˂lq��r'��i�B�J@�l�s[�5����`K��D�	a���Ӯw!\�8䮨��ekW���I|JHn��z��ea���4p���eqd���w&�r��VYW\�����[!�`�(i3%Ah�%4
>��XP����~��84Z�Ћ�l�TE�խ������S�0ů�x� ���rs�i�Vw�C�-��0#�tC%Q,!�;��
r7��(*h�Qf�kCH`=Th=mP��T�͌4s+�ny\D}��^��ٙ�D�s^E��S�Z鎬�������(���E�̱!\Z>�
6������+$��g��U-�e�v�W�G�[�^�������-the ���mh.�]����GC.�|���~��H��efm�0z�cUL���a��<mDrW�B��"���PB[<b�P�`<����B��٥P5���rs�i�H���N��C�X<� ���B��8�R�Z_.΄x�g��	��S8��UV��\Ƴ�r��Gh�Qf�\l{�"7�sa�vݝh�c�A�L'�1�d��{�ʬ�缆�YW)��͌4s+�ny �Ǧ�_@f���_t��R��XP���x���: �&�(E�{�ʬ�缆P �8�-�US�����U[�[B��$�����˔b�7D�EI����I�O��\�v�d�jFB��]͌4s+�ny]"Jׅ����d��.%Ah�%4
>��XP��Ȱ�^�7^/��1������p�V��O"�,�>E����\�v�VNub��pzl��a�Ʀ�|þM��a��zr,/'���Xw�j�7��r��&D�:f��:F�X?�g��U-�e�^.�@���e��0�U+�qbp@���K�Q�f�;�>)ʁ���f��Y�{'%sgeߪ�{ ^�x~�(vi�t�c,�q�T�\ ��-3zYIިuIF��^~�$�x�Wt!�`�(i3���+�J��Y�{'%s���䒼�7��Hn#���T�\ �͘�f��p�b�z'hۉ)���	4ˣF�n�5��cz^8������зq8�Ј'���Xw��fi~�'K�2��J���"�!ɺy���B���Ȇb�L���g�"�,�>E���]�!��	Ǹ�y85����@�`�8�Wǖg3ȓ8���/���fi~�'K�2��JHm����v�V�Nt�s$]�6����ޤg��c�n�5��cĭ#�?UM�!�`�(i3зq8�Ј'���Xw�j�7����o_��ü~���U��g��U-�e��)���UM`���R.OƋ.]$�t_-Z��T�\ ����Hq���F x>H�|�j���Iq��w�Ve�!8���\/Üy�a
�:�,�!��qƸ "g��z�WCp}��~Ϙ�g����P"X����G�"�|����.N����=��Ʒ����V�3��yɶ7s�9���o��S8����iY��"w�z��C���g��U-�e��)���UM`���R.���b\�#@[�I��Bg����P�ߪ��w��m�C�7���s��R��һY~����j��n�t�q�ٲ��+�J��Y�{'%sAX���	q���b\�#�y�Ya�I��g��U-�e��)���UM`���R.���b\�#�y�Ya�I��g��U-�e%uX���4N�|��Z�<kx8냞�!�`�(i3��Q]� _Fr�����WF!a�ޅNA��6D���K�Q�o{��:��(�[�*��Q]� _�rs�i��O3JT�!I�T�\ �͘�f��p�b�z'hۉ)���	4ˣF\d�RI��������yبw�ሑa7s�9���o7�B�J���o{��:�N�#�@j��{�`��Ҝye��B�o�\q�߈q	���S�[N��t�$Z���>�ߜ�J����^�_�J*�(��Z鎬������D��찔q_�pk����2%g�#0~��}�� л��@(�Ϯ(����%��yBD~"[
W���VYLl*w�{	�C�9Jn�+��Q]� _Fr���������0�@�U_� ��*ߵB`���!�`�(i3�!��@y��=�-Ǻ�:Nɲ`wl�����`�Ǔ3zӲ݌���������j��-�n`5�fK�Q2�+�Y�E�!Up-i�Cߋp{T���[�2ٛ�X�/R��:2QYeƈ�c�Z�~E�!Up-i�jK�o[���[�2ٛ�X�/R��:2QYeƈ�c�Z�~5�e`��9d��l����v�}���X�/R��rs�i�H���N��/Üy�a
���"X��[�p C;8;kѶ���� ZkIb!8!�`�(i3�d�٣�����6>�����ev.������f��gy:h+i
Z鎬����Ĺ#{��a'�<� \�Q�w���*��_?�v���Q]� _�:2QYeƈ�c�Z�~ݓ��E�I�Q�Тd�!�`�(i3�d�٣���,�JL���+ޡ)Ծ�/�n�*���?�#�6�fȯ�?
YT'���Xw�����C��'��/��࠮R:������V�6IWJE�r���秹��ч����=ў@'���Xwd�n]N�^ �7�}3��|�b�@a(􆿳���Qs��������=�8;�(�[�*!�`�(i3Ww�[h�q��!���\���Ȑ�'t��t�W�؏ 4�+�{_8�Y��M��)=໺(ӈ���x|}�|0�(�Y�MM��5��g�g�(�[�**�k�����\F�^�	E��߅�'e���婣	���U�dN�<@Iv�H�_��Q��b�z'hۉ)��!��|"/3�+��m\ƪ;���Q�0�=s�����[q�2�ߣ/s����.Y�[&���,�v����z��ˇ�h��ܙ�[-<�+�my$�N��YͲ�pzl��a��Ǯr!�`�(i3!�`�(i3�n`5�fK�Q2�+�Y��׎o�|���Y����!�`�(i3!�`�(i3�d�٣�����6>��i�X��*Z�!�`�(i3!�`�(i3�E����FZ鎬����Y�V��#qFL}��!�`�(i3!�`�(i3���+�J���q���U�pzl��a���gE��҂ϱ��[��Q�#<4^��n`5�fK�Q2�+�Y�kѶ���� k���3�F�-XX!i!�`�(i3�d�٣�����6>����9וP�;xB�_/�1!u7}:�E����FZ鎬����Y�V��#q胬<ċIX3�A���\�J2)V���+�J���q���U�pzl��a���gE��ҩ���;//M7$����n`5�fK�Q2�+�Y�kѶ���� k���3o=�<*��e���b��d�٣�����6>����9וP�;xB�_/]k�WM��q�E����FZ鎬����Y�V��#q�?�B��{k���3�z�Q�q���+�J���q���U�pzl��a�-{�*�;�Eo��K��]�q��n`5�fK�Q2�+�Y��׎o�|�8����|�M��5�!�`�(i3�d�٣�����6>��P��r��c� v?b���7;�Eo��K.�wK��� Z鎬����Y�V��#q{��>]#���)y(�O|�M��5����+�J���q���U�pzl��a�����;kn�P��l|�M��5��n`5�fK�Q2�+�Y�K=J��(��I(ީ���a41h���������d�٣���Ni�4�ڼ�t%>^��?�y��hL5ӥ����c^����
<ڑN���2�A��1��R�9*�eaA�|j?�d���&���>E��*�(��z�¿-ǂ,yߊ��b,�a������)�}�����T��.��W����t�.�!�8�}�\���;A<�SNp>�3������"h���ƅ5����5�`��N�W'�o����f7����e��x����#E`D���$G�	P��?[@S�CZ�~۵�q�#�p�	;�0�e�n�xdɨu �䆡X�dr�jf'��H������V���
���F:_ʣX`��_/��IC:GMG�2�3�A�E'����>E��*	Z�~(jm�7jl�N�Ar�/=�N�}���X	j�w~jiǎ[��S��_�:�R��h�4�b"����gE���Y(��	Q��H/!�Sy�+�z�}�-�%Q�a�4f�+�Z�{�b7�-�4T����	��,��<����r�k�,��~��U?'�����ٴ��{�G��ͫ������:[ۚܖ��`�[�	2�GF�&���#VW�GaAO'��7wT�,���P�&`bH$��>��L��$�I��i�j~>�Q.Ss�@�������-R�X��%�VB�=����R��(7�
��o��N⃟g��|"u8��d�w(�`��l4���/A� e8�~��f��Ԡ8�tF���)e���n�`�v�Q��7[32X|��h�ɑuϢ\�S&��)Q�����{1���	m���N����B�c���7zxs�ްs���	m���N����B :�Wd�O e8�~��<����B��B�BtQ���>Ft|�J �[�/��3Ɵ����s�3� BG
���L�}�J���2#x��X�	m���N����B��	�00�O�¶k��rH���G ^�����{ `�I7��$�ܫ �C_<qt�f�RUw����Q�h��@$˺/t��꫕qŧo��K�O�|/�3`�{�T}�j=�����dD]�Z��g��q���7���T��A��ˮ��
0'4\�A}��A�"�b���"v�����l������o+�@{fT�1�߽K}��׍���U�{'�$��'n�^0o����y�]֡�\�<7�X�e����yM��$��XP��Ȼ4�t=�j�.�/'��Y�
JHn��z�|=8�E<�l#�'�U(�M�z�v~S*��R��E����F�ҋX����@�ڗe'�c���9������5	��]�!��J�R�	۞h�G���4��'>]Z鎬�������(������ Z�U��c-a(􆿳�\�!��P�Q�$�k\_x���� �)b��X �<z�q�,+	�H��z���8�ϑ��[��勐�E�5orǟD�uiL${?���� �����Y~��`�J�,ˍ?]��IÙ=�H/��z��������m�!�`�(i3�b9����L�e�9%������1�;N�f�/H(TFGmrr��1��I�:!�`�(i3JHn��z�'>ftۿ�l#�'�U(�M�z��sّ"%4?e��#,Yx)�]�!��	Ǹ�y85����Z�m ��ߪ��w������4+�A!�N�By3��<Z鎬��������F!S�{r �<��z��}�Q2�+�Y�0=�!�hj�N�By3��<Z鎬�����R5�8g:�>j�5�i �<��z��}�Q2�+�Y��l-�%NvN�By3��<Z鎬�����c[��/�V�(^��<��z��}�Q2�+�Y�u:�)�r)Yl���#�]�!��荘�5V��ܤ�@�@y��v^�n����o�b?�����%a�E�IO����c�*c�r�w�����QV�i�6_چ�-�Z鎬������$��g,�k,^+a�@IE�U��w�B[��l����%T�� VU+I��V��k�'���z�����j.Z��$�sӢ(K�b	0\p c
N1z�H4l�I}}3M�C,����|#^�Vnֶ�����\P�O����X�e����M�:�'�R?�6��%]����	��鹾v�鳔��?�뭨�fv8���p�lő�4�`�+��t�Y�Ij���0E��@� ��L��Cÿζ]�HЦ����AS��M4m~�����c-�z��~��D:ǯ3�4���X�E��	�'�J���U�2Gޣסe� <���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9��~j5��Fo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+�S�AZL�0hs�A_	�K�o[��mU;լ^<���X�E���y=�$��]��	?{ʘ���d�kⲠ�([�߆4?d������X.S�����W�����C�"��0�����k�*�|*@l͓������yM��M��pAB����mݏ��A�)�u1Vp�߉n���R��oIZ�QCs">*���(�a��;�<�� ���2�jE?d�c���9��I����~uT`��R��*�)
m9��J�a$�Y FD�x%��t�oG7�=Ĺ��d��� U�����p
9}�Y�Ơ�C���"BC�I�1X����I�$�}�[���` t�:��������uO����(|u��W�s�ַ
���i�{��,>A�h�Y��6���]k�WM��qPs_*�GqW�w��fDf�z���H@�{���]K�I['�Ӹ��@?H2]�9e�a3 �*}# ����k�E��{i�¹!E��x�Q����V�/�h߲�������_����u�	"Ocbղ%�R��GN@����x�hn�B�l�2�T���)� �d8���l
߉�T&8�hbV�֎c�W�ƙb�;��5jjM�#M/Y�Z���$1&O�����i��;�~
���0�	+�����6(���j��h@S�@�]_LO;��Qz�#g�k���4+�A!�����;q�Y�f�ƥ�\����l�c���9��I����~uU�Ry�Ye��z��ic�s�yze�Zv�
!O:0��O�W�."��ђo�N������I8�h�N���&U2|5��/?Dc:���s�%�&�}!$ �7�]����z��z
��U4�i<���S)��{�R�$�V֩������;�j[����)�ޭ-�'h��Lc�Ո�D2��U4�it�|�AS�{�R�$�V�]�b��ގ��YWGզ86j�"Hs^�Z�cY�ZY3EZp��čb �F�gq��b�k������A��(aMq�P���ט�)Q���T�F�S~V]Ŧ���%��:7V�F�P�_�^���\�}�Z(Re]R:�8�����4����=�/!����'/�y=�$�̗�7�n�n3�#��L=6S�ʃ%�q�M�4*��G�^�I��rsM�T�J�b3Q���x�
FT��t����\�z���Q���J�R>�+Է̪h��|{�˕Qkgw��.�޹B$~s`�� �:Ft��m,UU����(M��&g;uA	�rx�́=5�ݳu��̒��Js�e�_��@��O@�*g����'�ȭ�n�h��� �[�:�5t�W�5=۟!��|�­�4h��K���B�q+�Ovf�?��$R�)�y�YWY�P�S��*Bo���+�竱����_�i(넃�<����v�/���d�h� v]&壁�ebÆ�����m���"�����.�)�r�S�<h�B*�2��ɞ��O֮�
V4�����}'� �>l+� ���L��ߨ�Vy��Lp�[��hV=������~�b"���$D@P�}��SY1�j�f?C�ms�~�E����	ݔ��m%۠Y�g�(��,|\��\�'�<�{M���)4��5傟�����O�{�"�a�<��ԧ:��� @P߬�1/ǆ������:n##���D�JN��D�k�e����zP�����@M��a�}r���U<�����[�(G��M��)��c�X`��_/���O֮�
�[�`7��pc �s��?���sF���(oW��;4i�Z"3n:�w���{찓�Ǹ����R�i&�V����Sv��rsM�T�J�b3Q��� #�`���q�X����B,'u��5rQ^5�yb��ޠ���U��%:��\�'ɬc��WN�ܹLh�l�|sd9i��mM�9W2�R���W��]�Jg����-0���+�Ax�`��v(��1��G�o�,·��4�w�j�a�N�>ˌ#�0�ݿ��A���p.Ey()v���v,�����e�xF����c�*�fsj`f�Q`!�K�UJ��:�Z~��X���RSr�Tʢp��Գ�AĘhTk���3j�;\E��ԄN���&U2����ǟ�|�~Ϋ�2
Ձi�ıν�7�]���&1f9m�҃�3���?�xB�_/�1!u7}:{�R�$�V��m5�@�uU� ��}n�8��D,^�d��d}'h����ć��mDm@<�9�X3�A���\�1��� ��9�Q��}�9��r45�`���R'�u)]��櫸�>ᛤ�f������9��|2Dm@<�9�X3�A���\���<&h ��9�Q�]k�WM��q�)0kcj1�kD�t�Sj̆��=�f�	�gȵ�]u(+֢���S,�D�c��Qԟ��
�A��R�j`D�����4m�1[�C�ߌ@ri��P��
o���;�Eo��K�p��h׬V�!+���}9��m;�n�i?3�(��J������i嶨��V����m�=�er߮�Ȗ�%T#�5��gE���؏{��ʝ�Y<6�B+�c%����â��[�J�e�C��1(�����d^_�Rꑽ,�I��a�|�j�h��K!/W��־�U��sp֟kh�W�f����C;��҇И|��,;���ͳI��â��E�❽�J!��8����|�M��5�М�\C�)1�ﻙ':]J�y�ZDU�.�Z�z�����b�y��־�U��sp֟kh�W�f����C;��҇И|��,�s0P_!��â��E���h�e�oM{r!:�k���3n-�Wfƍ�ѹ�OW����Ch@;���~q*��K!/W��־�U��sp֟kh�W�f����C;��҇И|��,N j�S�,���â��E���h�e=DmM�%k���3n-�Wfƍ����;y�O���[����0�%����M ���wi嶨��V����m�=�er߮�Ȗ�%T#�5��gE�����JԶ�.�I��$�w��<��D0פ�dV\p�W�\G���J�e�C��1(�����d^_�Rꑽ,�I����Si��i�rR�Z3�@�GݔO#�Z/��v
���M�wScp�)Z����(k���3]�b��ގig�q�M,@ri��PD���"��	���,��bJ�e�C��1(������˪Xk!�`�(i3��+!ݨ�k���3�˙	e
^�c���9��I����~uâ��[�J�e�C���Bm� ���M7$���b�Xrw��3�,�I��
���Ƀ@tl��(Ur��S��
	��-c��LU�L�����ج�~|�G��mO.�����R���oM{r!:�k���3�˙	e
^I�$�}�[���` t�:�yg��c|q!И|��,"��7Ch�m�;2Ϳɤ�櫸�>�����;kn�P��l|�M��5���U4�it�|�AS� U�����p��;�N&Pk���3�B�8���7�c���>��yС����І=�ra6yD�b �F�gqj�Ef��������FȮ�x]��n�ނ	��t?���`�n��U%aWp��.�替��+���<j��rbZƇ�P�X�;Qn("��94��On�AN�.���Ԃ�\�e��G����]�w9"x�g�Hz���m�W�w��fD} G��.��rb_6XC���d�k��h����S��s�(QY����|��[���d�kⲠ�([�߆4?d������?���+y��"nF^�{��s^��I�$nx떖ݏ��A�)�u1Vpйr�hr�W���M��pAB����mݏ��A��X� �:�.p�j(�KvMjm�f����qfb�B�l�2�����^t+��&���v��M��pAB����mݏ��A�8�2_�����Vy�G��M��pAB����mݏ��A��X� �:�6��ޡ+W�9u`�w��w�$�^�Q�[:Ҫqa���h�����,�ǰO8l5����u�z,�	��lx��Grkn��=�z#����2av����pJ�B����|��[���d�k���&=`+����t��w1�u.�����%Ὠ�p���\���`�+N���O��K��ݮ��a�=��d%�Z9 �VL�(\F2#���h�y
AHĂ_\R�)��<|k�݈�x�)NL	ٕ�����R�1��ԏ��R�)��<|k�݈�x�������yM4�"��2��s�5Xc�hbV�֎c�k�q��l�czD�k�$i{�7�<���qfb�B�l�2�e�St�F��6��ޡ+W�9u`�w��w�$�^�Q�[:Ҫq�b9�Y�y	{��g�p]?�d���&��n=:�Ed~z,�	��lx��Grkn��=�z#�c,?%�J���7#�w�O���<R�-�(Ktk��^�ѐ������m{J���F����h��
P�5��t-߱�~�0\��Ў�	;�1K��e�Igg�0k�,&��DZܤ�j&�+K���na��I�6��'�SS��gP�p=G�%�c�����c�,�[`��Z9`E1R�rF)���X�3c/��!�~^��/���f�;�>)�=e�ȩx��	�i��#�f�;�>)��)� �B��캧xӍ.��ew�T'+KK� ^���PG{��_�`��B�0w�]DWl$�`�]
���bI��2�}����2�����ǈݻ��y��H�W۞h�G���ڊ���$�R�<lͬ۞h�G����������I�&�`f��x�9�?�C<xWY�K��e�Igg�{��E0�DZܤ�j�]��	Hebm}3'\����2����I�}jI��C۞h�G���s�3����,�qm�c�,�[`�������(�;�H���oW�i��8t?�C<xWY�K��e�Igge�� �����DZܤ�j2t�ch���L�(�rY��'�SS��I?�KǶT�`NR���c�,�[`�-���u̳�rF)���X�3c/��!�p�O��{��f�;�>)ʋA���n_��	�i��#�f�;�>)�F'�J�Z~캧xӍ.�8(<���+KK� ^���PG{��_����S�]	=Q+����]
���bJz��.wrF)���X�3c/��!�L�q����f�;�>)��`�R �/�����
�]��2���ۖ��m�Υ,'���Xw�3φn �����m�Υ,'���Xw��a}���	�V�#!�c�=Ug?	��o+��Y(���8� l�O��R�(9�g#���)9�1v�1�9�$�� ��}�CU�+v�rs�i�H���N��F x>H�|�Wǖg3ȓ8���/�{=J���J��!�B�b]TF�����E]�:M�Z鎬�������(���^ �7�}3��|�b�@a(􆿳��Ri9�ꢅ�R*��\�R�&�-��)��\�<i�LE� R8�k��z-�%��u�	�c�4�b�E+8�D�q��27���{�ʬ�缆b0ؙ�02(�j�Z+�������x�dk/��+K��q;��x�gH��+�}&�~���i�x�^Z�wX������������4��&R��X�x��h��B̷��NfF�5.]��ȸs$f�<�JT_���F����7�<�
�dW���ֈ��tX���tl��(Ur�����398!��[
�p�F�Hj��]�3wN��JnZ�va�?F����M$]�6������o�t =�؈a������;R���M��j�l#��&R��X]TF�����x�dk/��ݾ-/̤�靤�}O�~���i�x`�ҧ��4�����[�dx �7�(��lj��
�j?�7r���g����,	S;&�+K���n;$�l��4�e���im�t�5���������J�Fbݙ�-M�O��~� ���K%����	x=:���{_8�Y��=�}�Vݨ��\9�oA�d��JXl'�&�P�2�PUг�|<Ѩ�f?�R��f�;�>)�E�zE�\?�([��}qn
V~$� +�,��݄����`�\���
�tf���!3@[�
 �ވ�*�'�a(􆿳�^~>��m�5ߧE4��J�1���k_���b_!2�͞nOYY�hg�N��Z�H�9 ���
�8��рa��N��*3M���*%C?*����l[j6�z���D���0�j�J�Ñ�����������g�R�"Ì�s��X�e�P�����`�B�I:׷�Fy�XZ@po��*���3m��U}�	��,�{�'�3�$ �#^�Vn���v_�"c�PƐt
�20)�_����*��Y~��`�J)����9	�(f���5�r*Iީ�4+�A!��X;p`�Z�^6Sծ��[�$���d~lr��[J�c�,�[`�u��s���6�ς�(�P�TEn1�♵~?R���v��|����q�is��+���Ã�E؀��<]c�,�[`��ᾮ$�YZ N��r*ً���N�c�,�[`�z�����?=7�}|��	���ˠ3� p�;H2��I�
�2���L�������XCk�8'��d+�����q9+t�}�c���nF�KD�Vr[?z%CS2b-M�O��~��s
!����p�>�q�M�4�%�VJ�F���˿1��;�H���oCO2��?'i��ċ�!-M�O��~��s
!��dʈ��Nf�ĭ�5���s�/����1?;��I:)��BZ��� 	1<�6�n�g]޳�;P���i)�/�1��P����^_曮�S��%[����;Ѩ�f?�R�����>q��A
��z(���7��R�۞h�G���h�T+]0���j���J�������ۧN�g�c�`�D�$0�Ʀ�|þM��
W� ���Pp��2�ĵ���Tzf��1�x�� p�;H2��I�
�2��f��U/(ۭ3�����Cߋp{T���[�2ټ�mˊ��ռ+���8�i@`:v�eQ~p�ܩv��Y� �(\�C����i�-M�O��~ӵG��b���_�1�J��]LB������%��v��DE8k ��Ck�8'��d+����'�^����&����1��⚺����jK�o[���[�2ټ�mˊ��դ�Hp9��Ԍ��Ǐ�c���w�I�7ݟ=�NM���ɛ�?ө�5ߧE4��rw�&�z<a��N� ��M�W8߸��S�Ȍ@�D�4��=R�.$�:��ż�����ӮvZ�A˸\MԂ�P���;>pRݴ�c"h�q�K�$d�A���g#�P|�<O����agz��-Cy�ݱ<s�� v}9��Ğ*��Eid_.lN�\���[C�}�{�6_����'��B�U�
6u��'KP���=� p�;H2��I�
�2�=�@)��۞h�G��0�=��l��j=/x9��g��ǻ�JLL?@J���q�D�*S���Ւ8����X��7L$]}á]�lEGV`2�'��B�U!�z@�!�~��Z2��u�>��{�����������g�R�"r�^K������О.�!H6F�� .�/'�b���' /�#nS#y����m�zЦ�+;4B�2��Ch`u����!��ٙ�D�s�U�V�Y\�J2)V���XR6�.���0:t�u��f�;�>)ʬ=߫>,I��3|�&�`ڱR̒�f�;�>)�(�W����<�Cr���X;p`�Ԍ��Ǐ�c���w�I�7~T� �}4�z�"x �n'�Wzp1��Xu������ 5#�3e�ά@�ș3�jn|��pՊhh�1-��\��Pc8;@#$Kb�i��Ӧ
J�RX�!��#��q�is���IX0F�M}���g4N�e���im��d��JXl'�&�P�2�PUг�|<Fw�1��o��xE�J�Iw�`�"c��k�nTK��|�!��G&)|{�ۚ�qSm�G۞h�G�9���n\�ӡ��A��h�T�z�Z�e�����1��X��WG ��ێoL�t���f��U/��s��U;4̽s�o�!��	x=:��f;[���x(�i��/Rh�x#�L_�(D{ͬ�y�4�����0��g��ǜ�-�A ���_��b�< q]����6/DX�3���.f{w��>���}{5���20{�(m�/i
�\ }Q'(�!��=k�Rm������ g�Q��Ȝxڣ9�$���>��o���Ώ<�?4Ck�8'��d+����}�{LFv(�c�,�[`��� U󤹼�j=/x9��c+
�i�l-�	�yH@�
@����=7�}|��	+�&i��V"s�ֵ�݄���'٥��gVا�˓#������N,=�c��m�>�c�Z�~J�1���۪	�}a�]�w%�oφ��<�6��'y�q�����2�,�B�����q�lj��
�jF�S� `�Cߋp{T���[�2�q+��=k�Rm������Κ?n���vF���M��J{�����qθ���7�W0#r�RN���6�Rh�HLN��tp�J��:�_�(�y�� ���f�hj�"��Ck�8'��d+�����m�jS��X��WG ���q�;���a*`�(o�l�V(��%J�bb��|k+Q�h'�Ȝxڣ9�$���>��o���ث#*�	���+����1��X��WG ���i��"u���Ȇb�L�($Z�u��΄x�g��	��S8�>���r8j�g����PTse��ͳ[a�<d��]��9��6�j��n	Y'F�0<gX����"�0S�l�%�z�J��3L�6(��dM�+���T�>���({")8�*IO��(������a@����L!�
�ݧ?���֭�Q�>^8�1�R@�e�c*o��ܔq_�pk���i��LKS�{�R�$�V��o{��:���m4��0�g�F}kQ1�8BW�R7���r_��m�q�;���a*`�(o�l�V(�ςMv!���xJ�1��슀.�[ ٓ��r_��m�o{��:�f0u�&�i"�ڬz����ɛ�?ө�5ߧE4��rw�&�z<a��N� ��M�W8߸��S�Ȍ��p|�
M
�q_�pk�����!Qr�g?	��o�dEr�+��#ȕ�B N��r*M`B�Ӑ�>�b��O�=7�}|��	c��N�o~#�ͫa��l�Y��QZ���$#z�*�
��Gk>��Mv!���x�o{��:���m4��0���f��J�a$�Y �c�Z�~����T��6\�4�@���(�?<n
V~$�,2�C�����d���Ą�Ĺ�,7�cL���	Ǹ�y85��֟��D�D���P�ħN�g�c�`�D�$0�Y"�g�YZ6��HHD�u��'J��l�o=��i֌]��	He$(�2�ft+�f�;�>)�;��e~]1bt�Z��P��3�Q#� :a�	�+4D@�K:+>%�C�5�ɇ����>�b��O������1�N�g�c�`k�J`�\A#�ͫa��l�Y��QZ���$#z�*�
��Gk>��Mv!���x7���.L��h�T�JDn ��aP�d�����a��R��q_�pk����2%g�p�X<m����a�z6�%�C�5�ɇ����>�b��O����Y5p��`Z"�A6"�ΝJ�Ut�\�W�{OEׁ��z\�Q��TXP�e�g�6�<+s'�^��������d�n5j�?�T�LW�_����V�&ݡ^����;q����}7�������\�2���.Z��'���:��KY�2Y��+rB�0j�䴑f��6�k�*x$6�ô���2�
�^��j"-M�O��~��c*o��ܔq_�pk��=��hX��9�{���J�sׯ�ɛ�?өW�{OEׁ��q�2��Kk:)���2��D+���4Y'�^����8BW�R7��� tN�y5�����$Hm�wS�$�����"��J�~�;�JCuym�Ut�\�W�{OEׁ��z\�Q��TXP�e�g�6�<+s�q9+t�}����d�n5j�?�T�LW�_����V�&ݡ^����;qf;[�����a�z6�%�C�5�ɇ����>�b��O��� @����ڲc�`\%����d�n5j�?�T�^'��s_ㆂ`Z"�A(sB.��Hf;[���Ĕ�.p�1��zB��݋����f��)�F��2p "BC�I�#�ͫa���n�e�[7�w�sB�ƛ��pP�����d�n5j�?�T�^'��s_ㆂ`Z"�A(sB.��Hf;[���Ĕ�.p�1��zB��݋����f��)�F��2p k��������Hp9���5ߧE4��p�-a�D͢fU�9��[b%Ɨ�k��"�՗�Cߋp{T���[�2�gu�}���<�f�;�>)�L��<z2���L�������]��	He\�\EǺ�Z=�du�([��}qn
V~$�s
!��$�ͽ�lF��-cL��)Ҩ�X,�v�x�GaO�]ڙ���_�z\�Q��TXP�e�g�6�<+s U�����p�zB��݋���>?���{��G�����{+��k�"r�q�;�Ӄ��g0?��7D�EI��o�D��%��v���c*o��ܔq_�pk����2%g����<-����R��n5j�?�T�LW�_��%3�o�:�p�-a�D͢fU�9�׏�����Mx(�i��/R�������a�U�ے
)I��%],=�$I�'���bp�7�ؓ��f��w�FZ�!>%/[�Z������-�1��~���סزN������<iwυ1�m;��g�0�ui�T�*�����j>Bj��rs�(�̴Y�{'%s�6F���y���'�'Q(Tse��ͳ[y*c@�e��'�^����ǆQV����QU�+J"�c�Z�~x(�i��/R�������a�U�ے
��]�U��!�`�(i3ZX�y�K�Ƹ.��v�!�`�(i3}S����inca߫r!�`�(i3P󯴈w1USQ.+��^!�`�(i37� ǚ�y��ɖ�~k�!�`�(i3Q@w�ӏ{?��5��!�`�(i3!�`�(i3&�{��x�l*�����l*�����l*�����l*�����$����!��Ƹ.��vΥ|�KyR��Q�!���!�`�(i3R���g����5�'.�!�`�(i3!�`�(i3�K��Oǘ����Fz�!�`�(i3 �|b�J�ll*�����l*�����l*�����l*�����l*�����tܑ��!�`�(i3�6Y^6ь�!�`�(i3Y��g�F�7!�`�(i3!�`�(i3!�`�(i3;Ax~?2����Fz�!�`�(i3��2}O�����:�2�����Vc2�����Vc2�����Vc2�����Vc���MooM!�`�(i3�K���I9��Ȇb�L��@]ˍ��JEgI�M�ĭ#�?UM�!�`�(i3;Ax~?2����Fz�!�`�(i3��2}O�����:�2�����Vc2�����Vc2�����Vc2�����Vc���MooM!�`�(i33��0��x���:T��Z=���KB�{�ʬ�缆(��۝} ;Ax~?2����Fz�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�4�!2d!�`�(i3!�`�(i3!�`�(i3G��0<]22�����Vc�R�
D~��2�����Vc�!n�'������Fz�!�`�(i3!�`�(i3Q@w�ӏ{���=��[cw�Yy5�����$Hm�wS�$�4�!2d!�`�(i3!�`�(i3!�`�(i3��%d9�^v�Ċ֩�*�yV�!�`�(i3;Ax~?2����Fz�!�`�(i3!�`�(i3M �̦�P�2�����Vc�I��+'2�����Vc2�����Vc���MooM!�`�(i3!�`�(i3!�`�(i3���|�(�����P��rʅ��a>A)��&�t5K����1��5��B4�����ӵZ#=D;r�R��xRGS��=[�#4�1L*��$#z�*,�c����GdN�8�g�;��|BT�=����_%D�-観�ݢ%]'\gWg�)���*�������'7�j�s륰�z*��['D�C�k�a�	�+4D@Gt�a�|���	x=:���{_8�Y��=�}�Vݨ��s��U;4���^a����HŹn�軑��r���/�ciJ�Kr���щ���ӮvZ��S)�3=7�}|��	��a-6�Da����b]
���b�-N�d�@/��r ��%�z�J��A`g.d�q_�pk��=��hX��9�{�������a�	�+4D@h�Qf��,2�C���s�Zs���U^v�Ċ֩�z��G�S٥P5���rs�i�Ǘ$� ��������-/J�����Ut�\�;|>r:w�|�sQ�:0 Y!܈��u@f�u\k-~ȋDa�vݝh�c�A�L'0i���crp/Üy�a
��-ײ��x���'RFtI��&� }iIB?�H�Nb�*Z鎬�������(���4p���eqq� ���+��'�����X��WG ��4ޓ���@�ȃ�ZK�9�e`M�x��h��B	���"�.\PM �%�s�~����gy Y!܈��u@f�u\�F�7A�c�}���Fo|k�Lb�"L?��ٶC$�-��]��9��6���ʵ���/�� �gj7�cL���	Ǹ�y85��֟��D�D���P�ħN�g�c�`�o<Z�L5���rEV��Ȇb�LH�cT֓O΄x�g��	��S8�>���r8j�g����P�A��i��ۉy�T�@.A�ov�rs�(�̴Y�{'%sAX���	q���x���:�M�C��Ut�\��ɺm7�{L.bC����s+N���D��N��c�7,�%����Q����ۉy�T�i��qol�h�Qf��5ߧE4��3t���=�4�04�jf�ɺm7�{�I���a5C�>��Ei�a�sir�@�A��I����!G�H�E U�Z��Tx�&ޓ�TpR0��ok%O�kai@`:v�eQ۞h�G�]t����qcR*E���&�Ut�\��F�R�M�ЯҞ{��6�.2�MWgX�����vs��P�<��^NEF/H�x]o/�� �T�1 Ҏ��7_]�4"m�u*w�Ac�}���Fo|k�Lbx(�i��/RŻ�&ǥ��a���F߸��S�Ȍ��"+VqS?�d���&�ق=�j��	�J�-D��`ʏgG�H���b��@|G�Y���J(i������`\5
�1��9��>F������>?���{��G�����k��k|�5J$s��(ko���Z��`펫���|=�
�^�^�{�`��Ҝ�h%�*f	�&�|��³��A((���ڔrcJ]�0���|mK�[�R?�6��'�|,kW�A��ˮ��V�rsSRąㄸKW�/�*��� [�	�z��7�b���W���H��rvXl�҂nǾ\�!f )[���Gs�������ܧe���5)Px
�B1CÂ������?k���[�ƭM��n�R�P�<��^N�q�is��g?	��o�dEr�+��#ȕ�B�������Ѩ�f?�R�g��j�([��}qn
V~$~�`������1��J�b�z'hۉ)��R�������T��6\�4�@���(�?<n
V~$_�)!c���~?R����I�
�2��.���-M�O��~��D�$0��;�H���opwI0����1��X��WG ���ɺm7�{L.bC����s+N���D��N��cߒ�ңui64ޓ���@\������fƑϥ�g7U�4<UQl��)I��%],=��m#�P��Y���E]9�3�c��?�)�||�-u��e��@�;�H���ow3Ԁ;M��1��X��WG ��>�7��=�1b�]`ݠ[�Di=&݇��I��R��B���m2 ��Qj;b��W���I��uP����by���1߽�\h5&���4���܂���:��KY׏�����Mrw�&�z<aSm�6��`4�04�jf��ܐ�}�S��/:+�e6j�"Hs�¨�h'�j��ͽ&�^������y�&D�H�B�*��QpĘ&�jW� ����!Qr�g?	��o`
��3�l�g�0�u���^a����HŹn�軑��r��4M̍����;�H���ow3Ԁ;M��1��X��WG ���>A�3�*��_?�v��g������>�wn��w��[#M���*����	���hKˀ�P��=��i!��ࡔ 4�UQ�}3doh�*��_?�v��q9+t�}Ż�&ǥ��a���F�LFC7�5$�)�vx�)��^�7=7�����bw��2V�RGS��=[��uܖ��m�el[�����N�9�?_��s�֙>�5�(2�q�is��g?	��o�dEr�+��#ȕ�B�������Ѩ�f?�R�g��j�([��}qn
V~$�UӇ��ɋ� ��X�D
CvK}D�؈a������h:h_Q\�=<�6>e��0�U+�qbp@�w�&1�|���yG~FsW��/dN�<@Iv��nt=:ྵp�!���Ct�w#��@t���3�l��d��JXl'�&�P�2�PUг�|<�D�$0�y�R�QY`�CgD�|A�$����@/��r �a�<d���u�q0O�*2t�ch���5�����Qa�	�+4D@i�a�sir>G���Mg"�jw�|�L�K�p��x��_�NH(�8��r��Ҧ\�02������\��4Z��՟��G�0��[��L�ΪA���Ǹ��St��h�T�JDn ��a������-M�O��~�4ޓ���@l��l��n��=���#P�j2E�?΃xI��o�8��9�.�`L��k�5��ng��	T�J�1��씑�:��KY���sm- _Y���@�}%@�`�4��h�3��'c�,�[`�t�)
W�k��
�!���i��ċ�!-M�O��~Ӿ9�d�L�<��lԻ5�q�2��Kk:)���2�u]9�#�I�X��WG ���9�d�L�� *�P���Ga��T�rs�(�̴Y�{'%s�6F���y�q� ���+�6e���mn
V~$�zR���b��C����:�ɡ�3��-e�y��FlJ^d�d��l�v+�öJ|-���{1�����ը�k:)���2�%��짐b��, �k��9�d�L��s"�k
�5��)�rbJ6�~��J�����ը�k:)���2��N�g�c�` e8�~����h:h_Q\M� �]vAy*ط��wng��	T�w�&1�|���yG~F�Y��WwOkd��l�\a���5C�tTi���׏�����M�q�)]Q�x��r_��m�b�P�LƑϥ�g7U\a���5C�o<Z�L5q�j�r�(�EoO�؁o��L��j\%�	k�N�L�K�p��qԭ(K�l���`y��+a?��J�~�;��1��Z��M���5^sh�Qf�΃xI��o�n���� [��ѮT��~��׺���d�����G��Ð�gxM��R,ng��	T�rw�&�z<a��r�����?0K,��=���*� о��PW��B9�[�c��)�-9�4r��g2�~������\��4Z��՟��G�0��[�q�)]Q�x��r_��m�i��"u���Ȇb�L��B bb���H��efm�0z�cUL���ޤ�Y5x���:����S�>��a-6�Da�b�P�L��c�{rS�b�8Z���%\��o���h�Me!d��q杳/��-0��3t���=�4�04�jfw�&1�|���yG~F�Y��WwOkd��l�\a���5Cc�}���Fo|k�LbJ�1���K���L���4�04�jfx(�i��/R�*�W�Ǹ!2�͞nOY�c����gp��T=7�����bw��2V��K粞ƿ�Ս���:��֭�Q�>^��(�S�����O��KJDn ��a��[�~ē�J$s��(ko���Z��'��s�"J�CJ+T �o��_�R�wَVݳA*{�;h/�0h�5eש�y�k�A�$����@/��r ��9[��meF<i�LE� R8�k��z-�%��u�N�^X�!ހ�����|E�g�������(ӈ��Z��&61�~���i�x�0mo��[0�ʂ�j�Ï��	�Li4"�	��z��R��Y"�g�YZ6��HHD�u"�T�B�Z�R*E���&�Ut�\�@�\����@���kJ���af�iβ�=&��]
���b���M��#l/����1��X��WG ��<a�`�&� �EoO�؁o��L��jDY޶8�1�Z3�z:�������n2\�,h������v�}�@(H�o��΄x�g��	��S8�>���r8j�g����PTse��ͳ[�%�z�J���h:h_Q\o�HT蔊�cٰ�Ž��v�}����6S ��x���'RFtx�W��L�rw�&�z<a��r����5ߧE4��p�-a�D͢fU�9�׏�����MFi��|ր���5V��	��yx�_uE���З�Df�H��3�L�N ��HE����P�M��J{�����qθ�)�A�������>�X���D�gZ�w&�d�I�_Lm����1Eu��P�6y�J����+���C��엫��RH[�3�s1����*�|v�|-J�g]���V�|�^���X���鰄;Sn;�i� �uC��1Vhs�`�1�O�u���(%�9QD�Pj�?n�3��ϓ�g�I�*MT�*��\���?��9)�F��Q�������D{+�>���3�G��( ,n/XE�{+;3&wӱ-���R�t����ʵ���$�Ƣ�/�J�w��|��1�29tX���ʵ���q���� $���{?tQ#���<0�U\�BJY��~���0����؈<�Ҧ+��U���J����+���C���ϝ�HX&ci�=hkrHo�??v�x�[a�в����n�q�^ƩW?�d���&���m!q��]�г9�=Q�|?�T�U)��4Ps_*�GqW�w��fD4^y@�c;T=0��:ƥ0����%���N�s��T��[C��ԭ��20`��WV�#aطR
�^0oߙ�(ml���d����=z��k�8]o/�� �T^��a�@�nx���:�owђN�~u*w�A�c����sL]~ц	U#�&|R�� r�l6��_.����q�is���IX0F�M��LV�!��o�½X5�g�0�u�R'cf����(-ЀU�D�� �����A�{2pn��gn|�P� &G�N�g�c�`l����d���=|%��v����a�z6�F�KD�Vr[?z%CS2b-M�O��~�Ѩ�f?�R�:��er?G��g��ǻ�J���G�&&�����@/��r ����z�/���:����嫋�T�@�.��KT��Ҕ�5Ɇܾ�]��	He$(�2�ft+�f�;�>)�;��e~]1bt�Z��P��3�Q#� :a�	�+4D@&����1�qSm�G۞h�G�e�ԑ\�#l/����1��X��WG ��Ѩ�f?�R�Ԍ��Ǐ�c���w�I�7['D�C�k�a�	�+4D@i�a�sir
>Rf�����v�}������Ja�vݝh�c�A�L'B��o彍/Üy�a
��ү�+ҋvE7�MW�+�Dd�,�alֶ5mL�#���+�9-�i"'���Xw�j�7����	=��h��h���LX��WG ���]�UQ��D�gZ�w{�R�$�V��o{��:���m4��0�g�F}kQ1��xȀ��D�[b%Ɨ�tl��(Ur,J��`�om�c�Z�~c�}���Fo|k�LbJ�1��슀.�[ ٓ��so�-c�,�[`����_�=7�}|��	��a-6�Dak��"�՗�Cߋp{T���[�2�S�o��VH� p�;H2��I�
�2�j�ڴ���a�	�+4D@vE7�MW]��9��6���ʵ������v�Z鎬�������(�����?�cc��L=X�� �-M�O��~�r�^�#v��.ȅ��J���B�:����}7�������\�2���.Z��'#P�j2E�?��˓#���l����d���=|%��v��3t���=�4�04�jfrw�&�z<a�4�ڈt׏�����MJ�1���۪	�}a��[�.K3�$�)�vx\n�ޱ��HF�V��r�Mrm�J��)g?	��o�G���k۞h�G�q���01` N��r*E����P�M��J{�����qθ����*j�"�A%o{?̊X����F��u��!}(`-Q�Xp�� ��~�y}i�#[<���5�p,[	jE�f�;�>)�w��9�������ф�ͪ��p�ϳNk���)�!,�!h3]1$��j�Ï��	�Li4"�	a�Xi��0�I���!2t�ch������N��۞h�G��6�mp�#��1��X��WG ������F��Cߋp{T���[�2�|�P� &G�N�g�c�`J��}0�^�s��R��$��_��cV׼�@��KT��Ҕy�R�QY�v��|���A�$����@/��r �,fc�i����r_��m�n��K����P��+7��]�����V磆�._�g��%X=����X�3���L=l���[��Z�q\�,h������v�}������Ja�vݝh�c�A�L'0i���crp/Üy�a
��ү�+ҋvE7�MW]��9��6�j��n	Y'F�0!�P.	ƒ�3^��h�Qf��lW��ڻw�;����<W�1�.����xȀ��D�[b%Ɨ��4�!���2�?̪���*��_?�v�#P�j2E�?�5ߧE4��zR���bѩ'�T<�ގ����r���Y6�Ei� ����23Y��P4,ժ �2�ι�^E��KT��Ҕ���{?tQ@.A�ov�rs�(�̴Y�{'%sAX���	q���x���:����S�>��a-6�Da��˓#��͔4�!���BC�x���}ip��`�rS�b�8Z���%\��oL�nU6�Mc�}���Fo|k�Lbx(�i��/RŻ�&ǥ��a���F�LFC7�5$�)�vx�s��:��=VU�簦~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢS����E@�gh1���Yh�\��q,f$�7Q0- ��Ck�4���_z�k�۸�y�uZoO�=���uc�A尋�N�N���aC�h�>1�|����ݱ�Ʀ�(a�&�����q��>��yܛ�	�����^�%k IÙ=�H�^�p"ORmHX���i�k�Zׇ	JHn��z��r9�3� �����Y~��`�J�,ˍ?]��IÙ=�Hz�n1:=��T.Ţh�S(k�E����F�ҋX����@�ڗe'Sծ��[�$N�By3��<Z鎬�����vl6m#�$
b��vr���(�
t��Y�{'%sgeߪ�{ ^�x~�(vi�t�c,�q�T�\ ���H�.WښBII��� ��P��s��{��E�EYZ/�矘��-n�̎�)6Opώ�,*y�#�45�{��	�FWJ�)T��Q]� _�rs�i��H���GR�>~qO�P��d��WMM
��,=��f��p�b�z'hۉ)q9L�Py4:��P��)��S�HZ鎬�������(���+��
&7����ҩؐz��6�����������=2��֕q1�r�5�Y�w����+��`s�;�E���nrm؊(�W���hnHN�~^;��?���z�����j.Z��$�sӢ(K�b	0\p c
N1z�H4l�I}}3M�C,����|#^�Vnֶ�����\P�O����X�e����M�:�'�R?�6��%]����	��鹾v�鳔��?�뭨�fv8���p�lő�4�`�+��t�Y�Ij���0E��@� ��L��Cÿζ]�HЦ����AS��M4m~�����c-�z��~��D:ǯ3�4���X�E��	�'�J���U�2Gޣסe� <���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9��~j5��Fo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+�S�AZL�0hs�A_	�K�o[��mU;լ^<���X�E������l��X�!�7φ��<�6�`
��3�l��èV;�jmT�#F�KD�Vr[?z%CS2b-M�O��~Ӹ�����& �^kM��K:D9����磱(f!�`�(i3!�`�(i3!�`�(i3�g/t��5����l/ǋq܃NQq�cl�j�)+�C�3�/3��
0<ȂD��^%O?[<��p�!�`�(i3�����L�	�=����k�\Dc}՟2[�����)i�f(7�p��'x��L��!�73I��o�
0��OA�t�U���j���J�r8�&=���������B�:_[�A��N�)��l�Gg�o�Ɵ����J�F�)-��.(M�
�p\,%�cy���7�!�`�(i3!�`�(i3�`�>'r�\%w%���Z(̼O=D���G��b�[6�'zT��2w�5����� ��=��hV���.�����_��D6��Ȁ`E�p����pd8����F���jbkAޚN��������~��ɳ���V]�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�$��@�/=e�ȩx���؛y+��:�"��m]�����q�c�'��D�o��Ow;t4t�f��(#����z�E��u1 )u!�`�(i3RN�]�5'�b1]�Q:~n�s~��20�OU�TG�eIw{������p�~����cж #���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g/t��5�e���!
�����_�X�z�51��2�nϵu��3�5�����g��ǻ�JhV���.�����_�uIB�+-8`E�p���$NDP�2��!�`�(i3!�`�(i3�it� B��~��ɳ�GV��)�m%@�`�4��t�o�ͱʺe��lf�F��e�m��R�km��K�~����c��C$Ԯx�!�`�(i3!�`�(i3!�`�(i3!�`�(i3nTxꅗ�~�K^M �ȸ��Q_K�W��m�/:��؛y+��:�"��s�n��c�'��D�%@�`�4����<!�`�(i3!�`�(i3!�`�(i3RN�]�5'y��$ŧ��=�qD�5��20�OU�O3���4�����p]��ܺ�C$Ԯx�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g/t��5�Y�n!�ƪU�\HU��\��J���nϵu��3�5����%@�`�4�$��T&����_$NDP�2��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��@֗�0
��� u�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�$��@�/Q��S����؛y+��:�"��*��\��g!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3RN�]�5'�b1]�Q:~n�s~��20�OU�۾�\Ը����p�~����c�;Ym���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g/t��5�e���!
�����_�X�z�51��2��K�G�5�������Oam�hV���.�����_����˸�`E�p���������2�!�`�(i3!�`�(i3�it� B��~��ɳ�GV��)�m�7Wx� Pa�t�o�ͱʺe��lf�);��<�O�R�km��K�~����c�<�?���!�`�(i3!�`�(i3!�`�(i3!�`�(i3nTxꅗ�~�K^M �ȸ��Q_K�W��s�x�62�؛y+��:�"��6���BI�c�'��D��7Wx� Pa���<!�`�(i3!�`�(i3!�`�(i3RN�]�5'y��$ŧ��=�qD�5��20�OU�J�(BJ�����p]��ܺ<�?���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g/t��5�Y�n!�ƪU�\HU��\��J����K�G�5����7Wx� Pa$��T&����_������2�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��@֗�0
�;���7���LFC7�5$�)�vx�،��Y�C�e�W�0��D�����	X%+I�$�l'�7��ܓ��;TL���n�3���j��!�Lc�TH������7��!j�L-vc�,�[`�_k����ۧ� #چ��+,	����sCݗ[��ޭ�l?��n�5j��i͠Z��)2��dh_��tCv�*<"��� ^�x~�(vi�t�c,�q����Uh1�� �:&��L&fL0