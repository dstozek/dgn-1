��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t����j�X�8�����$4L�������}g7l�� *��I������,0�z8O� ��t'�O��!y}_���C���cC&��BB�m����_�2rI~�K0�HR3=�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K��un�ZOF���_i����T�3��aO�����V���n,R�L���>���
�&c�Qrg!����x�
�%{2�c���'է��7�u��ursf!���͢^�sܻ���@�3���	�����/E�u�T��I�1Q�A��DqH(X1��~^�ۙ�����{���?�k�]d��0��kc���8�N��D}�.؝��7
�h	aڍ��*�:�����Kw�� w��ГJZ��1Bb<p�-��X���I;3cd�N�������H�4۔Cn�-����>�'�����;p���J���Vb���&P4x��V6d$�?Ϳ��ҕ�����ůP3ru��@.v�)i'��W��j^6������]N�T.I�=r-҈ג y;oZ�V�?\J*�����ޑ;���������*���v���=q��W��XvkK4|�6� '���C����{=�a؈w��F���VV�w׻�����,����ѢӟaU�Izy�k���?�J`���0��Mzᑙ��Qb�^z.�gO`��	�6�]s1�@i�}�=�����aئ�Ͳ��A=��Rn#~���@�n�*���W,���ͷ}Ŋ�.�E�:�,1��4`.��rO4�MK>>����Ԛ��#iȒ�$v��ǽ�G���wla��������u��$�θ���ĸ�-�v%�&�Pr�-���D�qhˇ�JM�ڽ�y��
���;��	 �Lr��8�z�M���À���f���@����Аx*v�%`���I��L��<Y�x�(7D���_��a�$ &Ҫ���jgR��_C�Ԧ��ОS�D�y��D���+,�2�x��O 3Y�*Z�G�x��`�@���jVMM.F������&Н2�4�e���Ht)��6�au/#�����4���3���_Ey<����`�M������ ��"#���f�h�2�p�5'u�����Nh<*�gY��T�Y�+='�Ԙߜ����*�����'8yʖG�S�Lri�&�$٢w)�h��,�5~��Ti���n�	�	ju��'�{��|Q��z�^�H]8��	]*��0z ��e�-0�k;��������W2��'`\Jx�z� �-"���9��x*LiaD�p���U2�t�!�O�4s���2���ǲ9��瘆yJ3�+b��YrC�01'ʥ��y�#�9��J�|ќ0W���M�W��4\�q�$�[�i�������|yk��b�"G�6ASz����ױ��8+v�H�'>�n��#b�(NO�׈��Ԣ�/�7���َ�Q�3���b4�N�$��9 @7��Tޢ�6�;�֯��j	����R^Φ��{��/��K���������N(�k1�sk�-Å�IM�T��ʝ�����%
��O�Y��ż}��SA�a�*���.�,��χӓB��$b���=�]��U�{޸������rR��ryO�Zͧkx:�������ʥa�=�m`���S�V��2������.1��j�f��w7����Y�2$�)G��9����i��E���b%��;v8aŗ��3j�m��X]��@�B����	�i�y��h�u�ɩsd�������^f�K�u��a:�z�'b�ء|sU G/Z�m��?�>B��;����9�jE���H����y�W���L^M�
�`;��5��5&c;5�]���2|j�p�R*���t�Uf�,�@���	�ݒ
�@$Sb�4WY�#���v#��ݶ����W�CoHp0�W��T��|����¸t�A3�7����??�t��&�P�'�p`�d�:�X2����6�;���& ��iI���0o�|H��l&+��)n+R�A:�Cy\��(��l�m�g� a��^�u��F%[����X�����kN _�~��\�=�*
� T�y�P���d�9� ��O	�58~�=���[Jf=�H_a�ϥUb��ڟ�"k>J����� �)�y��Z�#�0��ƵE������*��S1a� �X�\��_b�C��v�EGke4@�{���ӱy��?����8v��_��i�P	���'���Ęj~n��i�^��[��v��%!��^[0l2�60��݇�K�s�΄.W� \�bpܩ�M���e y	&\0�!*�jh@����d�W6��5��g�`yhk]�-i!�<	���,��.���6�zj���6~�	r1�
����#����<�Sڿ��1A�y?7�� �k�j"y�&(�b�I;�^�;��G�h�қa*����l� _rƵ�-���s F�r;β�	o�=FX!�g��հZ�H���l���]!}��Vkܕ��ң�V����[�,�7
��K$�u�l���m�|� 
k+s��1�6�`C\�?��|Ko��ܹ��j�+D<Z���	�G�a�n�pE������b�
`ܾ�7����㹁�=>eN�qi���.�T��R��Qږ�/@��e����j��0�˸uAҍ]2�/���.�(�.g��by�'?|L5[=��O�����k�RV�u�
���e����V�R�����K��g��g#����
tL�\��o'��-��ؙ���iԪ�C�PnW1=U�մ�{�i��5�R�ݴ$�B
�؜���F�G#�/p{0�wQw:����� 5�e��Q���f�4Q�a��c"K�R�l�#V~ڏ�U�`�0���B��Myx��Y^�FO��8���a~2oj^ljw�WG>&�{=�Ǉy��+�o�Q&�ԣ5)�4��1�A��ۜ����Z�p���ɾ��[�+�vR=�34"񞊀�$*#�~�b
�.�`��;z]��Y��$��7k`+-��9 ������e�D�u��1W��~w�[����d��wt�Ϯ�Ь���dΦV��P�k�;ˇ/l\�ғxR���+��]@/��)�ɠ������(!��iO��e^��;�4�y�ʌ7���ca���M��?>�V3�>gW�ԧF�jh/ˍ�
�\�*�lTA�wxt��l�jiG+�$¤LRn�[$��xt��K&��S0���K=�*x<Bt��p�J���.6T2K{W1.���a��Dٟ������F�Q.Z3�hU�I�J�Δg��@�Ѡa�`P�{	!�
�݂ Xt������.��L`Y��ֺ��k�L�9�}� ������8ɢꏤaj�*ӊeN�u	G��A�sc�S�Cˬ�a;:!����e�C�J�"��&<�[#8�c�E~z��_WV�F������hf'��ts�����`R��	������7[p@��ջ�"kv ����B���Q�z��pl���3�ѩU}�&]~�}>�"�`+a� ��|��"�z�e/��8���PM�]�bGO��n �zcRI q�.��+_�5� 
�vn���Ds�椰O�~�';�c��J0�\�	�5��v�m>L��Co�&-߶w��n�銑�U����N�wu	�"(��Ճc6ks=YBk��l2zU�a�h��1b��w[Ժ�=o�܂(\ST�|�|�-�'��r\����=}%���1Zұ�s�'ҿ`1!��F4�V�jEBn��0Ch(*��ԢS`N���Y@�	�b�Qgg������
������?�d���x����q���d'�5�>� i���V�쳐AB��`C�im���(�f���-a�EY�QzЮ��gʏ�_�7����V�\W_��"�'m;�Xm�LVU$�-L���� ���m����ѩ�������yOt��a:�/�+���B��"��彫ّC��j'9��(�)(ݲ"z�Y����WE1�L��ws����,壘��Ka5>q����Wްd�ȏG�lj���Z���i�^�� M���8�Z�h]�co���IA��r���4U�8ї�= F�Jz������t�L<B���*τ������,}�<���-�wa�CN?�eO �H��^8\��d�m�T�����f:�u�I�KF�����ѴƎ�I�R����3 �Nn���*�=έ�ꩍ|�������nד�*��.g&S�GV�%���0, l���u�Tm�-yvd;������-Q��'�����H;���d�:)�9!_�@s�:E"H�Ш=�/׀�qV5l�́��H��TS��_��1"=�SF-�[���5ț�RK��1�SG��[���F����-��+��%��2�65\�j��NN����.�v��[�Jk
8bP�6:.s1�Fz�h�s�)���|��F�m�K<53t��_�d�L��=�9
ZU�y:6m[��f�u�5�P�?�{��m�* \���d#�}#�qRA[�A+�!����d� ��(�@��.~	�XL����nQ��NwB�^h=��b��g�bN~�E$�s�nw�KR_�Dh������4����u}ٴ"!e�S뼼'7n���%)���'���X G�fq���;x5"���=�c��}�J���y:3�/�l�'=��4.�jS-�KORd����R�4�s�drʘע��b!��@i�~������K^�}T�Ul��6pP� q�+1rЍ��O�� ��#���tmߘt���^44?�\M��[������4C�}H�'y�kI|KӸ���>S/�R�:Q�
n4ob��}������u�Nj^��K��h_������y��b�-�s�$]`7�z�q�
WE���Xl��|;*�KUiꬡ0)���3eHxSq��n��Tv�N�W���2o���B0��DJ�:��n)_�M�.l��/�߄|��?i�߫��)�]�lg`V�+�e��VV�+�d�QZZ��y��	4����R%Q��/"
���@��Y�U�={�����}�D���0��Q��?�ïJ��P�ԧ��0�lN��.���	���=Ӻ�yݬ��JP���bH�y��C��Hd�� �\�TM�Y,;`��^# ݿAtQ�7X��aO�%ՅlM[;�����^���kT�QX^X��O��8��U@�0a�ab��nr���� ��g��AG�L�����.���I�_7j|��	����p��D�X��/���;���y�<��p����ǚk�W~������(�YP��	ށ�9Y-�a��jtx�ڑӖ��Xm�eb���nT�W-�G#��jDa�W;�5 |� k�Rۮ�u,q�UG=� -~;D0ZŵKP���8���t:�_�����ZMh|U�C���6�9M������5\�OZ��F<��U�gB!<X�ݰ|O<�7���jƻ;���%FX��I�F1�����
ǖ�}�����p���Ǡ�9�u��y[���E�a�N��k
k������F��^�p �;�-���[!����P�L����!��}a���E�Zġ�zH�')yW�c@A���%����+���5�IOO��gŸ��n����m��4��*�+h^����-+����DGb�WI�J���7��uXi"�cLT�-OV�R+1o|��0������'U�h�)��L��3�}1���:�y1IOh�o��.�Su���C��XBB|��u;^�ϸ��xR%c�d�-J���@t�nM�n��P�P۾]hA���hHI��{%��7R�V[���r'���FS��E�?��6'I<��fJ�1-x|����<����I�����u<�A=��F��K��h�[&W�\w>��h���D�ژ V�^�s7�7T�?���w��ыL��\�!��QÏ�T�$Z�`��n�ܞ3�/1��.�����*;~j���^b��&z�co�7q�������pM*p�u�Ӹ�-�n+�}�<��D�\4�Dp�/��3*#TF-a��塟x��r=�C>�b�QHM�_(+��-�/L5R�M�Kѯ{�@�ET9�T$8C-v45����5i�<)>ʌs���Hh�؞:�����DlX�����mDM�l͞��f�6�9����O�@kE+�kg�F�&����a�O߃�#���~o:p�ښ�j��ѩ�K�&�*�� �\�p�J�fN��k�5����{�Nx�ߴ�a�����"�
Ӳ�wL'�5��b���9���M�'����c���)z��郿둶<'����pIH�@0~�@d���u?�8?X�)�r>�ǳ~N�G�R9h��A�a��E�k�ߟ3���i!6(t��ڙ�EID��_~��-
��+�ߞo�y���ݕ5��n��?%!�^v����5�duV��^���-e�/M/����-�v!p�C��z�9q.���4�ð���z��f���iD�	���^� L�5���!�ϵ����~����r^U��m��뮸�⳴��u��%��|�N��}��#2���ڀ��`Ɯx�H��u��!�����5D�E�4��o���9������k���� U�e�����㡚��G<H��%��d��C�9��&
���ff��¯䞷h���������6�A����QT����s�GAZ��5G�FPzs]���ɠFo�Ɠ�%�A؋3�
u�n������yR��J;�Ap�6�!��vP�6p��Ǔ�Z�P���,����놺32(+.���m�"<PYP�s*R}hb��p�W=�a�{Y��OK�\؎"�1r�L,�c�v9YO��=G:-�,�����)��(���6Ң:O��q-�jD(�GI?Ak�rG����DL�]x�8��V����+�T  ��,L�of�5`��0��fr��Z�+�n��t�Ͽ~��̓q��L���le�J�U��s0�ɉ0+f�����s�^��$ܪ)�K��J�[f�fA���V/E����$5|xwe�=f�3�10*{$�3
zp��$���``��%p��3+-!�I뛅�+� �7cŃݮ/��a-��CoЙXO�1q�� z�9�uz�E=��%b�u���p�$x����q����
�<��Q�͝���P]G4@��e��Я}#��D�3Cѵ��<���s(�|�e��w���� S���KSW>���s]��?5��gMNF)�P��F��LF_N�)�\�O Ve�,����>ݐ��9ѶX��J�V�|��h�x1�S�kf������.E@���ւNl�=]]�s�.�d`��	DbA�_[ִ� ��ӕ�c�s� �9�J+Y<K���U�r�Sq�5@y�$�J��9��[��R� ���rߏ;br�g��������@0̔�r�5<�8�T��
�`Ti�F3�&m|C�r	��$NNq25=�G�ƱN$���t?CW0%��\�F���^^��-��u��q�$U����/ɜ��n�e��x<�K0I=$@K"E�,�N��y+�`��.f;|~�hѩ�
�v�K��Yalz����ڞ�X���^~���]�Q���3L��na]B���@�f��8|A�K�w�3AZE2��Em���,�@�Qql�kPOkM �w��-h�V!t��Ӟ,}`��~�)�ud�2m�p��5���I�@Ǥ]�	�X:RYbaa�i���,�ɟG���d�HO@��:�{��g�ahܾ�����W�A(	�r���w$�J�� �i(���u]����/�d|ҽ��j'ET���N���ĉ�tO3^�	mP�*Xp�]�z��)��ȊU�0+r��V�(_����w<
��$�w�w�B���$lǫBA�8�a���y��'v���ᒌ	�QR��*�Q�(���G^�Zd<0+-��Ss�!#�;��O2yW��Ë�場ݰ����AYbt� Y}	���O�����Mw'���>����0f�
���z��;�b���\{�g����M��$�Mp�)�H��}��*h�H��ԟ2�}�n�,E�euP� ,cK0�?�!4wV7:}l  C������z��1�S�r��lv�sxs@�
�Hz��|@:i���Ω�B�Q�N�� ���R�M^8Rqׇͅ�:���\R�)����0	�1+�5<���hFrG��ߺ�3ִ8PK].�:�� �� �xhT�НnJMo��^0�!���Wg���e`�-Փ�W��U�U5*�.g%�6)��.8y�qi!\���(�ޭ�=��:\�:*^���T�������e�i@7<��?��A�y.cA��za�;.���L��ގLɤoa;�F]��|wr�i�:�D4��{5���4]Vj`�@'q�}�E��&�(�i:���D�K�J�2��&[4=L��#y�+i��!�i�J��(�f���� �X����&�ϔ�s���'C~sS2�S���o��uQ5q�sl&�}
Ϥב�O�3�Pd�n^�,M�!m\��"�Iia�����:wY�$���@��8��R<U����g��T�-�C�S�ub3,ҹ~z���P��F�؆/�$S�y9�Y��^���>5]�ts�9�t�p=�2�So�nDTg�0�R�u(��PH7�"�]��!'o� �_#?��$:��L�F1��Ejň=5D��-P�w�@(�T���5���m�&��'�z}��<I��CUn6H���iE�כ��h�����*����?�N�K�s6{S���!P�M�q��m���oZ����l<���|��
�J�7�J���G�E4�/��K�b�kM���J��-0��Hf
Y��Bv H�ƕ�����:�Oͼ�D{�󷸃#Q��
�Z4�|$�r����[�1#g���Uv�zD��c�1��d�"��H���Ӳ�G���NR��Ϗ
����T ���ҿڶGs�	/j��dw�d�o@	�� p�=��D�e+�Yh`^�0P�H
o��7�?F�5�N���	F��=�?�s��Q�p�URC��u���:���Q�ws`��m! ��o���U6vb�����:���j�C�Q�Rft��e��2��7����b�k�.�!�g�VY�"zx*U�+v��$^h5��œ��A�(>��F�۶�-X��!��)!]�
_��Qp��vh1Ծ�|t��Y���R�D��Ċ<�	E����K�X.lSp����
�yP<��6m�_��Ǝa� y�]�Ӓ���`�$�D#� 5O�F����|��D��c��eG��N���s�Lu ���`�����H�_Й(Ҧ4D�/L8������S�w()��£�pX(�Ry|.^/6۪�1� �]� ��CoڬR�xO��[��ggڡk>�[_G�ʂY���=Y�Ta��sP� ��m��b_/$s0�<dq%#�4���u&[��'m`ѳ���c�)f�V#5J7v�bc9�(����Y�-��.�0C=����ۄ�܎h�,�	�@�g9�Mӑ��#Z�*g�,��,;�ϿU:���քHGt�=��LÑ#M��}�^s�?�u�(c���!x��9a({���\������x��Y���������Q�84(��
�̹�˙Ȳ�hG¸�Ci�s���R)X��ꚏĊ$d��+a����y+�[��5Ԫ{Iܓ�N�!�|�1���/�<G� �-���!��w�Cº��>��g��1�=Ǧ��Hf��}���Iˁ��X�OK��x�$��m��Eġь�T��ki]t�r��/��#0�Ѿ�s:FN��k"���"����Y��\��8QP�A&�F�#���1�"0+�:*��1�5�{��ZL�M���Ee8#w\�5�����Qҭ.��zh��c�ʔ����@:GY6��U�lA�4����蛺_)�"����I�?�1�%��U���>"���{�C������6`�h���������o�\Ϊ��2UZ�H�-3ŵl� ��w"A�
�V�"�V�������F�A"Ag�}��Hb�.�*\�b�-�ǜ��(V�-��i�v�l\Ҋ�n
<��D�܎P�r2C�j����ֵ8\��Β@ ��e���D���=�T���G���
}�Ͷu��hc3��WQ�<�&�0�k�b���e�Z�ߨ�=J V�0l�=U�X���Q�6������l��_6<�)uH�6��ך�d�"����� ���NL��E�x˂mYJ��D
*߼�b�e^���ڗ���*W����);I����̾9 U��u��#Xd3��)�@kU�d�˱T�G�<�n�))�dzݗ'�<‏�:��W|�<�;u�KOa����K�����V��A$ ��H8#�����f�	B�aE�L+ӎ~<����h�b<栞�y?3ؚ9�[ܠ"Y�K����P\}�-}��>�#���y�ڤ�$cV��1�!8o�,m)z����g�����o�c�8%(! ��I�����@��8j����9��K�Kw��ļW�e��^"��o�0�r��;�^�ť�3C�JN��.���x;����^�����9���i�M��O��2�s]��7I9|�?VG��J�5���n���	R����9f��h���z|�z�vN�2s6�\�ѝ�����UX��\I�8s,mY\a1p��RUjsݫ�0�X)p	�HAY�/d]rq����f7�D��V]70C��@Gc43��if�o�	C�'haHL*R#�� b��N��ӔK�ﲐ����"l�J��5��� Hv?�ſ�M�J�I���k�#/ۆ
�K����Zn�5E�ӡǶ
�:��Y�b*</�@��pD�>"��K��J�~6�jg)�	b��&
�^S��[٣�Yt�DT:���h�&�*�0��f~����dܹT�O���ǋ�Q���:ˈG>D6$�����D�@;�,h�
��!�3ƻ�R�hR�4�u� L��a�8�͡fO&y��}���T1ʷ[����;�<�%�;\�5�7d�qMg���H,QWL����6M?��B_��	��+O��0�"0c7:x���sN ��vH���A��c�^���!F^&��#�f��݉��`Qm��� F�D��6!���kT�|�N�)�l�Y�݇_��M~����}	�m(<��#"�$��Ά$`>��`&�܁�,�<>G��s�ø�����FHm�$�~�W��hb�~fm���R,0�k1��/(G�YOz�s/��֫I.(������n#%<%��R��E�)ϒw�٥�~:C�ȓR^>h��bd�ݸ|�p��=]ve���XRvuyN�Ќ�/v�JI�5:�x�5