��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-
Ү��p7Ȩ-Mw �)��\y���{�z�ox�!P���b6�')Ri��_�
h������a�;5B5Y+� �i7�sp>1�*_��h_�
h�'ʯv!	��;5B5Y+�T�����N1�*_��h_�
h�Su�X���;5B5Y+�0�T��:1�*_��h_�
h��!n�x*4�^ֻ����XP���3�Tt
�w�}of�O��p�k����\�U�q��&�'n�^0oO,�����5����`K:���K�n̙z7��(�Ԕ��~��'n�^0o���{����I��'�S����cܙ��u�X����W�,���Op�ե[CF���y7�5����`K:���K�no*��\MI2#H:�d�TpubMpIÙ=�H�{	�� =�R���c&;�/��V��WB��	K�U�&��9�Sca�&'�'n�^0o6��U�x���5����`K:���K�n̙z7��(+�}�Ҳxh�믳��"5� �S��Z ��d���%�a�A��CN�vs����L ��xQ7��y��Vu��s$y�4�Dg2^��I��'�S����c��2gF����Z8{�):;5B5Y+� �i7�sp>1�*_��hjOhi��ȫfc<�R{X���w��|��kVU_�E�I��'�7w����w��Z8{�):��W0i��^g��F����%�a�A��CN�`ѽ�N��}:�E)�F����@��zL͊�q��K��e�m��0nZo�j���
,H+�Ӂb�9�f��W0i��^�A�hA�@O1�*_��hjOhi��ap���
)��;�}�u��s$y�4�Dg2^��I��'�S����c��2gF�����ͧ���Tq{�f��a�P9b����%�a���錜c��=�
>��$0�"��	֧�ǌo�9񶺸��_���׿k[Ai����@0���u��s$y�@�~T�@��5����`K:���K�n�Z(J,��*|��:\��^ֻ����XP���3�Tt
�w�Ocm�r�?���0�i_@#�8u��s$y�6��ܡ�.�5����`K������*|��:\�+��CY�E2�e�.�
11�*_��h�����T��u�{��2.��p��3�̘*T	6�'n�^0o _xB�I��'�!f_\eN�g	M@�����W0i��^�A�hA�@O1�*_��hjOhi���Fϴ��hۃ�T���|��N�p9:O�I��'�S����c��2gF���^�iq��;5B5Y+�.��h��u>1�*_��hjOhi��U_�8��oْ�h�R��|�����j����I��'�7w����w®^�iq����W0i��^O��bvq���%�a�A��CN�`ѽ�N��)&%�����!����q�'n�^0o{?�@�I��'�!f_\eN���Sq�`�2�������Ż?�N�`eg��Ocm�r܉�k�־/R7U��(�"5� �S��;��� ��%�a�A��CN�`ѽ�N�����C�H�^ֻ����XP����`eg��Ocm�r��(�Mm]�_T��d�P�?��{	Q�L�`Ȝ0nZo�j�B�!jEx2U	���:���Op�ե[CF���y7�5����`K:���K�n�Z(J,��&��C�<A�fBN.):�
IÙ=�H����������׿k[H�1�?$J��X��[�"5� �S���
y����%�a���錜c���B��hM�;�v��u��s$y��	o��I�5����`K:���K�n�Z(J,���L��Lv��̍�59�\��\�v�w#<r^��|�5����`K��m���L��Lv�Zή;X���u��s$y�6��ܡ�.�5����`K�������L��Lv�Zή;X���u��s$y��	o��I�5����`K:���K�n�Z(J,��&��C�<A��=�X��h�'n�^0o@�~T�@��5����`K��m��&��C�<A�������92��|�����j����I��'�7w����w�ޔ(�w��_T��d�P�?��{	p�Uh�9h�5����`K:���K�n�Z(J,���L��Lv��=�X��h�'n�^0oP�Q��([W�5����`K��m���L��Lv�������92��|�����j����I��'�7w����w���Sq�`�_T��d�P�?��{	f��Y ;��͌4s+�ny�Gz�SQbʛʇ_�^��Ů&�Bq{�f��aƨ:bN�t�~[[z�'KlJ�D�5���L�gp1�*_��h�����T ���c��_��١9�G~��ڹ 	�"5� �S���
y����%�a�A��CNשY�w�ߒf�[ۻƆ��YGQe�.��Op�ե[t�v�N�͌4s+�ny�Gz�SQb����=�s�A"&Gu�RA�uS���|��N�p9:O�I��'�S����c�W�n=?Bv(�J��)��)r��>�f֧�ǌo�9�3*]��@���͞�^�x�����tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM�f<�,=K�F~�?|�[_	E���=�[4�l6�Pr"?�8��	º��%�	�r�)�u&ȵ����Z�(��׉󾶓:��,�w$�z(����Ig`i�'n�^0o����y�]�v�'�
Δ^ֻ����XP���"Ru2:#g����3ê�C����\�v��62,۲�XȨ�@PPKȶ�/�l��Y ���#�w�3�0���F$��P�{��H��[��d����;aY���H�q�4^���	���嵓P�?��{	Q$�fB9��9?_��=Y��_�0z�cUL�jk./<�6���{�c���
È!�Z鎬�������(������yԵ�Z�n��[��{_8�Y���˂lq���"B�� �ƽ]dN�4JHn��z�:�&���Ϯ� л��=����Ҽ�pC�\[�*n�#U?x8�Q�l��t�KS�#�͂G�ƥ+E;5B5Y+�+�����E �d�n0�+h5�u���Ͻ�Zı\��4�޸�b}� �y��~�f�'n�^0oڀB��:��	aQ�� xS4�q��~�<��p�=�������_x�} ���>���{�|��	y��~�f�'n�^0o�C�~��j�4�aY��`ս�B���dV<4����;{ۤ�&�TF�jK�P��r,�e3F���);�%�N�YE�WzL͊�q���,Na�G��geEq�l���j��I�:iZ�Q����*df("(���	����5:ղg���sq{�f��aƑ�nt�� �<�6�Q=����W�j�ZϚ�ڊ=�B"��jk�$����v7�'^�J�_-�_3#ڸZ鎬������Eu���7P��T�<��z��}�Q2�+�Y��\�6�(�_3#ڸZ鎬����N��q���$�7P��T�<��z��}�Q2�+�Y���3�Mo��v�~������]�!���<:���u�����~��|��].��'���Xw[���YD��Ig`i�ҋX����@�ڗe'��osq��|��].��'���XwMb�+u�b;b�4�L��_3#ڸZ鎬�����ǥ{��{��L�9�r.p�B*�2���u���d�ӿ�>��f]��A�5d�HР�{��}�D�T�٥��T� �73w�tU`f�g_3#ڸZ鎬�������(���kk�ȥ�S�}���G��Yʬ`�f��`y���̬���	p��[�6ߝ��{2l���^���@�B��Es���.P������͞N	���m�]|Y27� ���֕tx!����^�i����(�
t��Y�{'%s2�ew�S����c����.q�B�Yj1� P���������(�M�D�bó=��!��L����犷��r��\Uo"S�%X�hZ�0�`�ò��Ҡ��Nr�3P���WT�j
�I��w��,�"��ȝ�Qؚ\���Rz/��C_�#��2���TC�<򶁥��9�dMbZ鎬�����aC8��-���^��.�m$�֔ ��[�M$�,WʿL�TD���9�,�w�-�
֩����gs&�~ס&���#�{�0;�}�^��w
��G�Z�4{���a��l��0xCv���p�5��\l��,\ަ�It�M:��2�w$�z(����Ig`i�'n�^0o����y�]VŤ3+���;ۂ��IÙ=�H�<��S3�q�4^���	���嵓P�?��{	�<��S3ϣɻz��wSx�lޞ��rs�i���H��	/���{�|��	k
�R����d�٣��c�A�L'd��������Cҷ��e�ˇ�h����2�[Qnk��XH�U����f3��^ֻ����XP��ȣ��hg©Z���� G����Da��������/�%疷���-���^��woT�c�\�=�1p��'n�^0o!��0ך��$��o��}M��`�ܜFS҈�l���K���q�[�W���^ֻ����XP����5�2���d\��7f�%�'�����-���^<fGc�� BD�Ai`�}���O����{�c�%l� f�HIÙ=�H�����*m�iT����(�a��������Pk��)X�b���,S;���~V_��(PyZ9���{�c�%l� f�HIÙ=�HE�]�L����r��=W�6�-z!-x�n����WF�B�[#�S;���~V�Ծ�ʰg���sq{�f��aƑ�nt�� �<�6�Q=����W�j�ZϚ�ڊ=�B"��j���=��s��{`�s�# ;����Ig`i�ҋX����@�ڗe'ٜ�U�n~q_3#ڸZ鎬�����R5�8g:��⿣:�d��{l�f|�ό���.�;,o��1��č�Y���S�)37J*u)T{6T'��OG��_3#ڸZ鎬������E�^��L�����~��|��].��'���Xw�����2��7P��T�<��z��}�Q2�+�Y�wZ K�Ϋ�v�~������]�!��f�%p k�yd�A����W�+���z�ҋX����@�ڗe'����vA=8ܞ�}��z��eU�e�����'��E ]ohWt�_a��7��;� ��Jzv4�܉-`�6�Ԧ*��>���w%e���{l�f|��rs�i��=29��a��>�\Ԍ�m��H�^��"X��[�`�L�i�e�	q�X�ZQ:���U]�Jg����-c �ЄW:c��;�&����\��z�+e0���0��h�B�����2f�ƶ`��:BY����^�i����(�
t��Y�{'%s2�ew�S����c����.q�B�Yj1� P�������^���N�Cp!!v*!��u���d�Ӵ���)�jj���|}��i��{��s��N�}oT���zV8c.K����Ig`i7G#+��Q2�+�Y�6��GJf��誆�J �$y�;R�����3���Ig`i7G#+��Q2�+�Y�m��|�Wgak��s<Gd�oaL�!�����z�	:�WT�j
�I��w��,���|HH9M\��e���S��k�U��i��16��t3$��z�9���x���Y)�x{0xCv���pSFh��Q;�im���M:��2�w$�z(���!��ZB	��5�HT�����E��<K����Z;��1й=�$Q�r�q�4^��ɪ�nj��L�aG�>!�!���{�c��*�^��\�V��D�.����E��
Z����\f���<UA�>��d��G�ƥ+EǇg[����ĉ��0 ��[�W����nj��Lv� )�j���{�c�J81�%��}؇ld�Cp&Zc��g}Ю�0s�# ;���!��ZB��,�Ӏ(�ٜ�U�n~qbS�xǠ�j�đ4��B�⿣:�d���φc���zT������!��ZB�hiY�����3�Mo����v·�t<���JY�mݶ��h���X ���@Wk-ɢ�����t{h���X �<�h<}�N��osq���n℄o.�h��8�I���d��I��v�R��$k�R�������K6��%����_$W{���`��:BY����^�i�����m�q���z�n��9�n,]Q�yfT�9������h4c뻖*����u��z�	:�h���R���M%��3+�7�����L~΄gO�3f��*��������[�/�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@��<��W��k�۸�y�uZoO�=������;6��ȐTo����'p�@�k�U��ʧ�V���,\ަ�It�i$�$[���ɾ�;ۂ��IÙ=�Hb�����K2�:�5q{�f��a��4�6�tڬF
��[lD�����.(��"5� �S:Zot�{> ���{�c���
È!�Z鎬�������(������˚�9��9?_��=Y��_�0z�cULL�֗ul?�T�\ �͘�f��p�b�z'hۉ)r�k��)愥���ޤ7��;ۂ��IÙ=�H�42_�'
�7eUshl~�Kϯˏ�K�������ܭ�'��:�^��8�m�\�=�1p��'n�^0o!��0ך��$��o��}M��`�ܜFS҈�l���K���qb�%Y�w��;5B5Y+� �i7�sp> �d�n0�����9X�O� �VI�:iZ�Q,��\D�ш���g������E��Vib�%Y�w��;5B5Y+�T�����N �d�n0ϙ�K4`����j��I�:iZ�Q�K�3X"��6�!��w.�4iI��d����|	q.�q{�f��aƩr*�^�	�<�6�Q=S�W�$E5<4����;{?^�Z��μ�P,Uw��ZmM��j+���0%ђ ��zL͊�q��J4����(���H�Q���12\p�G�iAL��K�~����.j�,�3*���Xf�.�7P��T�<��z��}�Q2�+�Y�ٜ�U�n~q_3#ڸZ鎬������	�$Y�ł�u9j1�f<��z��}�Q2�+�Y�塂
Z,�_3#ڸZ鎬�������En;,b}����[v��{l�f|�ό���.�0=�!�hj���Ig`i�ҋX����@�ڗe'�Q;�m���|��].��'���Xw�m�l"ƣ���Ig`i�ҋX����;�ƀ�'͚���6�S:$���H{R<��z��}�Q2�+�Y�����vA=8ܞ�}��z��eU�e�����'��E ]ohWt�_a��7��;� ��Jzv4�܉-`�6�a��x�jT%q�#�<��z��}�0z�cUL���gM�6�!�u��އ�e���3a(􆿳��b�zx����� �*u�,-6�41�e�LZ\^ �@'�ZX8�5}7���_UVp
MMo�����!Au�U�l�+mA�g9�țH�WT�j
�I��w��,c�A�L'�f?S��##�'�\�ge��T�\ ��@ #JڃC����a;�/8'�L
�2�Ot�ky����<04�ΟO��n4#��Ԕjݭ#����P��:@n��9�n��(�
t�ژq���U�� �`%$��#��� ����hѓؤ���3���Ig`i7G#+��Q2�+�Y����P���k��s<Gd�oaL�!����lY��qq/8k>6s����]�!��$��lW�d&� ��JL��{� 9]�����>P�2-i_���F���/�� �*	��q`g��Iٞ�߹��S��|�s;�'�o����f^��%e���=<�HITH���cCV�uq��T�6s��bk��d��w���=F�����R��GwF�|���&��,h ��o����j\�|��܈�7�ol1A]VI��	}����ā"�z���J�v �xU�M���l�������.Z�.^�![���8�v}�1�C��Ÿ��at�������@���>^
*��?O��&Y��V��m��z���d��N�s��U��=5��6�0O�@�(>v5�=V+��+AF\�ۡ�7���+9�0�eh�G,�LТ��-�{2W�ke� KB�~�.l8��� �5i��$ۏ���I[�ܯ)�}�����T��.��W����x�]�V���_�;�W����Y3[v�8�>P�2-i_aߌdW���p���q=Őn�C�K��x�mbѿ'l��$���wT΁>����+/beGIUa):nX�Y�L�r� 
����7���w��c�Q(�u�8�Ix�,bσ4�^�ϷW�(��$�$:�so�5��m�w趤ې�3❡�<�W����N>4�~)5�(���{�eV���C�T��,Ny��j�_�>P�2-i_�d�Wz|�D]��h�	�I���(���Yޭ�A�,�����5�����:�kw�x��P�ɗ��A�,�����;ɾ2�� r��4��(`��`w��ANw+���A�,�[5[��6��N*�x��`����%���Z�q�N�hY!=��8R��(7�
��o��N⃟g��|"u�Y�CP+MdPuʟ�1K�G��ئ�#X���55���F�� e8�~�� ��!~�2O�R�<�Uh�*�bh���d��fs�B�d�K����H�S��x���Z�1�s�;�2B��y,��6��ƙ>�_O�S��x���� �>���y�9�d/Ѹ���� l�ߎ�����-�ku��?�b��M'���Xw�j�7������>�u��+�v�|B���x}�E�C �۾�0A�!S�UE^����Cҷ��eYVf�c��<&��s�z�A���f�}���G�QO�K�E׼�\�v��<��>ّR�vC\��S����c����.q�B����GϤ4�s1�&X~�u��8
� �^��%Y�g���"R�ݪ��֌??^*��7$��Q,�!Y�]���KXͯ��<�ݢ���|B���x}�W�\s��t��J=;��5����`K��$+~�%�Ћ�l�Ta��k�����)^G�<�zL͊�q��VR8Z�ڝO}�K�=�����S��7SYT�Rs[:��YZy� VU+I���=�e-]���Y�p+�@{fT��+��z9�f�G��bu��MT�	;�HIIż�\�v��:Y��z�i#@���%&E����T��;�Ӣ����L��1�gi�q���U��� j� ��/%ѕ�KW��]�!��5��E0�ؚx�ǂ}���X�7G#+��Q2�+�Yɷn����b��8�hNq��Z鎬�������(���R��F�D�g��U-�e��,�R�ܤ�@�@y��}�6�����\P+�}��A�"�|aR�A>T<�jo��f�\#+��SВ#]k�Z' ��뎆Q��18_��i#@���%&���$�O�C�n�6o7V�1����]�!��	Ǹ�y85��^�	 �wa(􆿳�tP"7��%e��0�U+�qbp@�%c�f�g��fSg�MEZ鎬����d+����NG� ��j�ҋX����L$�����/'٥��gV�HZJ��ݢ�{l�f|��:2QYeƈ�=�<�^�-��1�R4�:��*'���Xw�����C����۫�����tK���I��w��,���|HH9M\��e���S��X�l���4�j�����U��_ڊk�窝ה�����oP�^�u�SC2R+d�8Dѕ�O	ڰC\�6@���c�Y{�^�T�YP���sA��$���Xq֧�ǌo�9��~��l��g�'�� ��뎆Q�P�?��{	�i��X@�}�K�
�4l�v �?���	�sq��17G#+�ǟ
��|�6|�+�� VU+I�O��v|2&�d�;o력�oԉ�hҌO���orǟD�ui�+��V����"1{"��\�v�<A��s]��5D܅���'n�^0o%�vZ���M����$�l#�'�s��P{����zɥԶ��{�,�I'���Xwd�n]Nِ����_H;a(􆿳�e�&���6!6�ymCoZ鎬��������F!SJ3��Y�z�Z鎬������E�^��Lk�np�h��]�!��V�,�q^���O��U!�Z鎬����b;g굈�Cde��0���q���U�,؆Q��4�<��z��}�Q2�+�Y�]���P�a1@IE�U��w�B[��lQ�$�k\_x���� ���CZ�cQj�d�䏡e4�1H$�DZ� C�C�.�.ܟ��		�bt��&����d�٣�����6>��s��k'?	��-�2���=Y��_�0z�cUL��]��~	�}���G�>򵘆m���g��U-�eu�,���$�����3���-I'��~����oHq�p���\c�/峞�<@��=Y��_Q2�+�Yɼ,I_E�6b���������Ig`iZ鎬����Y�V��#q�s科Df?���Ќ��=Y��_Q2�+�Y� �r�54�W���"��[B�����'���Xwa'�<� \Y�F#Q	p����3�]�!��	Ǹ�y85��~�g���` �f�N�g��U-�e5��e6²���[�OR��K�c Sx�lޞ�ό���.���K�Q��0�a�����k�]�!���1����m���[�O��
z��>Sx�lޞ�ό���.���K�Q$Z̐/[���Ig`iZ鎬����Y�V��#qe+��4��F�+����j�ﻋ-���C�M��N��e��>O������{5Ø�=Y��_Q2�+�Y�7.YL�7��d��IMf���9���q���U�pzl��a�@�=�)E8��E��1Z鎬����Y�V��#qV ,�6 <?�k��]�!��	Ǹ�y85��_3�i�GT�#��+�������(��� ��d,1��5C̘�=Y��_Q2�+�Y�"��+����Pr���mSx�lޞ��rs�i�LZLø�ʞRW����Z��T�\ ���|.�TӏE^&�T��z�f}�tL�]�!���1����m��w����9=W�玞���K��pzl��a������	���嵓'��֔�����>^�2�����Vc2�����VcREBR�hHr�A��5�V�����w)К��g: k��2�����Vc2�����Vc)���f���T��+{�0��WQ��I��L��%��v��h"&;�(�	�����M-я&��x�T.�_m��{�R�$�V֦���ȫ_V9�GKP�2�����VcREBR�hHr�<;�yr���1�vt��9�GKP�2�����Vc����]��pP׳�A"*�A
�7�$G���s��DX@^w
��#��+��n0�)�^?�d���&�������ײ��lP>���g��
�٧�\�T�q�>�YŇ=�er߮���^��oF�v�മ#F� �gO;\z�lE��p&p�Wq�1~ԭ�@�Pd	���~)�iI�
���1vs����L ��xQ7v!:Ӽ��t��ж�﹈�iǇg[������u'K���%�ϗ�w�/EI���āsp֟kh�R�4>A�}0"�`�ҏ h���X �) �c�%���(M���9����,�ǰ��ZA����}���������J���6s�,�=����+'u��ɛ��`���u�{���Eny�\�fl�3Ys纁#g�k��B���({`C�GD�d���k�窝הْl��]�B/��v
���+�K=�Jᬉ>:&�h���X �7w����w�Z�7G�}m�0�|U�.h�#nn?l×n
9�.��_��C��N�'�m���1�R�M�&H���١9�G�29a���Q\f���<Uȫfc<�Rm�"2�/EI���āsp֟kh�R�4>A�}0"�`�ҏ h���X �) �c�%���(M���9����,�ǰr�
\��;AO.�� ڽ��
�1%9��4��aA�=����+'u��ɛ��`���u�{���Eny�\�E�tF ��4����>�/�����t�f�7���G�x�l��1i�t�U	
�̔�}͑!/0�D��nj��LAi�����̷�X�Zx���b��]���;��d;��f��2R!�u��އ,),U2�CM��G�j���&"���vIh�e�B>l�2��!f_\eN��n�s�۱�*U*�������S,�D�c��QԶ;�Ӣ����a����vE��HT��W��ϼ^vc@[�_zβr��H9����>�/���kt�5=�=��	E��/�*�>��"�$-���`~[[z�'K�8�t��O�����ҏ��Z�������,n�*����IY��j���[orǟD�uiM���	�fl�Dߠ˨�R+d�8Dѕ��e�������*|��:\�0�|U�.h�#nn?l×n
9�.��_��C��N�'�m���1�R�M�&H���١9�G�29a���Q\f���<U�|H��(@�	��A�v��GݔO#�Z/��v
����vH�fIA�����N��v�R�ZU r�_]٣�2e�tV��	��y}1Z��2W�\�?Z��<�I���P4T��ʬ�[GO>��-G�r�6���`ѽ�N��)&%������%I�@A��~�����d�r�T���t�f�7���G�x�l��1i�t�U	
�̔�}͑!/0�D��nj��L��㴀@�^-�2`s_�]מG�u��t��?��CG��>�\Ԍ\$⨹�2H�Q�i���IK��m�F"&[�Z�{����m���L��Lv���l��;�4~���;A����z��%c�f�g���V��\_G($�y�&@�sZ��|�+��?�d���&���8$E���|��ˏ����_ V�z/~�a��L�Ɲ���S����c��2gF���b�V�"�;��|B�Dv�ەRu�8Ҕ-RH�y��-^7]fn�c՝_�\�Zr�D�c��Q� ��c�M��B5���^�Z;��1��B��hM��<�U��B���y��Ţ�Fnź	P6���:l��,����-l��e��+׵�d\v��s�#%�ދ�����nj��LH�1�?$J����&4	�/��NO�l����m�=�er߮�1Dg�Ŭ�!��ZB.�,��G�)aޫ<�:$d�c����,�n����_ V_/J��6�- ��,"J�Yǹ���O��<RʉGO>��-G�r�6���`ѽ�N��)&%�����Y
�6OX���#g�k��(1�G#?Fpe��*�Ǡ{u:K�����t�f�7���G�x�l��1i�t�U	
�̔�}͑!/0�D��nj��L��㴀@Op�K��l/u���!�P���sA�el$gS��:���K�ne�rE�*o.:���p�+~����f�[ۻƆeu��<̮Z;��1��h/��8Δ�=D�0T�/EI���āsp֟kh�R�4>A�}0"�`�ҏ h���X �) �c�%���(M���9����,�ǰ.�A���d*�<`#˟׾��.I"�UJ%`�}l����c)9+�홹���ޠĀ�=����+'u��ɛ��`���u�{� u�WA�=�lH_���U�C��k:w�������l�\�B��xC8ՃA�[�Y����AW$��,\ަ�It}�0�.�,l/u���!�'���UV��H M��� B�!jEx2��M!{S����b��]���;��d;��f��2R!�u��އ,),U2�CM��G�j���&"���vIh�e�B>l�2��!f_\eN��y�,r҂8�/��NO�l����m�=�er߮�1Dg�Ŭ�!��ZB.�,��G�)aޫ<�:$d�c���4�C�>\h������l�\�B��xC8�FvO���a�������.I"�O.n<~�)���IJ�.i��ܰY�̄��&|ù1,k�T���P��?�d���&��Y��/ �s�����Yǹ����u�}Ԝx�k�窝הْl��]�B/��v
���+�K=�Jᬉ>:&�h���X �7w����w�ޔ(�w��_·x������@�Pd	���~)�iI�
���1vs����L ��xQ7v!:Ӽ��t��ж�﹈�iǇg[����I�u��ZnH������*U*�������S,�D�c��QԶ;�Ӣ����a����vE��HT��W��ϼ^vc@[�_zβr�)V��B�1�f�Q�:���[$�n8~�"C����w�X�.B�s(dA�+�홹���ޠĀ�=����+'u��ɛ��`���u�{��2.��p��I��8�>�;��|B^E?2W���mM�~��+�1Dg�Ŭ�ɛXL�ڠ-RH�y��-^7]fn�c՝_�\�Zr�D�c��Q� ��c�M��B5���^�Z;��1��3��JS�M�~��t�kE	
�̔�}9MpW~�b�B�GQ1{��S����c܊/��8muS���dWk[�W*e/
Y��g�'�鶴���;� �gO;\(��OX7|�df\��'�1�/��NO�l����m�=�er߮�1Dg�Ŭ�!��ZB.�,��G�)aޫ<�:$d�c����)�f}Q��?V���qq��u
��yrY��B��L����d\��)c��S+�홹���ޠĀ�=����+'u��ɛ��`���u�{��C�*����JwYu�%��?�d���&��Y��/ \��)c��S+�홹�����Y��j���[orǟD�uiM���	�fl�Dߠ˨�R+d�8Dѕ��e�������&��C�<A�s�4B��ǆ��J�`�Ӽ\���L>�vHUHN�ʯ$�4UBQ�/�*���jš���:Q�l�H M��� :|'4�e�2��J�h{oZjF������(f���i�t�U)����SO+���
0ͺ���^lONp��q��-�8qTmI(x;��|B�#��f륖9׃�&�I��Yǹ����~{yj�C�V�4�Xape��*�Ǡ{u:K��px�$��řynK*�%v:���K�n�Z(J,���L��Lv�
a�o��@^���\�}C�V�4�Xape��*�Ǡ{u:K�����t�f�7���G�x�l��1i�t�U	
�̔�}͑!/0�D��nj��L��㴀@�L�gp0�|U�.h�#nn?l×n
9�.��_��C��N�'�m���1�R�M�&H���١9�G�29a���Q\f���<U�+Q
O��	�w���)O�*U*�������S,�D�c��QԶ;�Ӣ����a����vE��HT��W��ϼ^vc@[�_zβrrZ�0m�\���O�̧�	9`�����yrY��BQ�ߝM��'��<I!Rғչ:���K�n�Z(J,��%Q��&����F� ²Pt���^��r���%���8����F��C�՚$9�˴y�?����ׂw�.�G3�E�3��.����]�w9"x�g�Hz�N�1�� ��2�����Vc2�����Vc��Y7�к�C4�M���Al��H��>��\��g: k��2�����Vc2�����Vc�cRq>h�^N��l�5�/
Y���	}�@��4�wMh�` �f�N;��|B* ^���x�>n��L�XN��0��X��wu�w�2�y�����b^�N`���H*�����ƶ0h�5e�J�qC����\���fb~*��s�;��hS& ��} �ZqzO���Cð��T�º�������H1�q9+t�}2Z�<�����/�ciJ��
�5�������h��)�kǇ<�<���Hn
V~$2f�*�)����3�s��{��㐜��xQ�n
V~$d]��>����Y2j���]��TM���K�+EC��t2��9:���K�n̙z7��(��u��V�n�%�z�J��������L���_u-'٥��gV��"L?���<6�<�>���Y�y��2�嫋�T���Hp9��x(�i��/R�P�HS|�4�04�jfJ�1����ݾ-/�uu��ڿ$�)�vxe�zA��;��|B���.���� �2�����Vc2�����Vcl��w&� ���!��K
�M;y����&2�@�2�����Vc2�����Vcv�iL�Dqy�e=��bƓ:H���Y�pQ;�im���M:��2�29a���Q��nj��L�Ă��������,g�k0������ܸ �gO;\.��R������M:��2��!�_b�Ȥ�J#��9 ��.]����hl' ��ߝr����|��T;)��LrCQ�i�r�ӯ#7�k:���I$��T�ķ��QԉM!����sh���X �;"U��wF�v��n�y�b�\D�Ix1W�fB)����N�9!��9���9�GKP�2�����Vc2�����Vc��Y7��$�^��ۉ�å�^1��&�,���Fu)n2�����Vc2�����Vc2�����Vcꑈ����hfWs���@�!Ss�7"�0�0�h��#g�k����W�세��w#�1�b�z'hۉ)��R����=WS
���q9+t�}@[�_zβr#^:ͣ[7�k��
,X���^�%ʌ&&yR7|=����+'u�ֻ��K���Z��ᗺb���M�I��օzUo�Ӧ,\ަ�It}�0�.�,�W7��c�r )$"��-�Z;��1С0�U�}�:^�+�J�h���X ��S�������~�;����ɝ\�!2A�C�=�.��*�{�ԅ-�1Dg�Ŭ�!��ZB.�,��G�)��r�n������T%��h���X ���0�a��[�����ɕ2��Ȅ&N�/.�B/#M!����sh���X ��U�~��N���\ב�wI�6g4�xhp���D�{�B?���L]٣�2e�tV��	��y���p8��RM"���Y��ݣ��2�oesĘ>��*�����Ɲ_�\�Zr��<E�Y�*eu��<�Ǉg[���ȉ���S��(�2���s�;1?�[F�sp֟kh�5�o�|D?�J� 	Z�ģ�{ucN%9�%�Y�`��3*!���E|�P�t��)OA�����Nh���R�ީ�����M��j�Q���h���X �y�������h��l|�ϖA�#�l�B�u+��h���X �{Ē���o�ߍF���!��ZBǉ��'�V�N�\A3
b�kr�^�0:���n�b���ڧ����h����0��}.*#�}�J��X��+�d�q�^!�`�(i3����~j^�q�����f-��9�K�1�!���:���K�n���SYƒc������С".��H�	��	!�`�(i3<��Q��\��jT�):1�#��Н�3G�J�pD�4�n�7$��Q,�!Y�]���߼u��u��s���'~�!�`�(i30��w?�h��(Z+�<Vo�eopREU���'�WkjNY��##�'7[8�i��JU��j5�2�����Vc2�����Vc2�����Vc�m7���e,�����?ݤ�RD:9�Y��f���Fu)n2�����Vc2�����Vc2�����VcϷ��6D��}|�R�R��G0�6f׿����q�>�Y�}>�x�t4�փZ���0�wU��=�R�̙z7��(��N*�u�[
�}3��*���1������1n`�{à X( �H^��t�x�n�[�O��_���wg�W���'hN��;�Ż}����[v��$/��>���4w�g�P_��'�!��o�V��?"��Ho�d�	r������oE��cFl����h4c��+��#�v���`4�E%h���R�ނ6�l�yŶ��띚<�74���o�[U$m�a>�JU��j5�2�����Vcv�iL�D��_�̵<��� �\�遦��Fu)n2�����Vc2�����Vc����0+C70;*��/c�W�BƲNu/T��� N��r*����_�{`u���3������7�\�&(�B�s�%��v��B�R���>_B�`�� ���-''�����.�,��G�)a�d�X.9�X��WG ��Z�e��0�뷿ʒ������3�so�*s�Ԃj�ߝE r ��E-�%J�1���۪	�}a�]�w%�oφ��<�6�'�-�Ss�kD�It	U��@�!Ss�7"�0�0�h��#g�k���V��M|8Es��pUo��l��n�4��0����?�d���&���ʷ�JZ��!��,S/� d�Rfi*=����+'u�ֻ��K���Z�וzj7i�j�70;*��\��!��>�j�s�-�(��K�M���u|�M��mW�e�(�68	�I/��\]�3�� �f���c�>�����f2g�d�1c�o���$[ ��TSG�7��$Z̐/[�'eD�֟�e��LU�rw�&�z<aSm�6��`4�04�jf��ܐ�}�S��/:+�e6j�"Hs(�R�A(�
Rygv�_��7���8�i�H�\� N��r*d�*qT����Y1k��z%a>*<UB3) �c�%�<���Hn
V~$��0�a���I��q'q�����N��ӱ�WX`u���3�U�'�]�0�Ú�On��m:�yI��^]�Q�I�^$D���q!�E��q0t:O�G+̈́�J�����3�s��{�����4y��ijX��WG ���:u� ���a��xK�0�������w_��{��e��˴SI���x(�i��/Rh�x#�L_�(D{ͬ�y�4����F����%2B�܎���UpG��|�'ݍժ�\�Ȧ���0+CjB����C�G9<=k�Rm���]�!
��!��~���=7�}|��	�7���:���
��c�Z�~�ȴ��A�v�i�a����w��ΊB>���<���Hn
V~$�$�@L�Xd������ݾ-/�uu��ڿ׏�����M��ܐ�}���e�x�f
�[q�_X=����3�spu[���7�\��}���.�����_�G.�
��Y�y��29�R?3S�j�;�J�/�y����[�O�E�B�f	�l�;�:��(��l⺬sw'%wy��$ŧ��K�A�2G��k-�^uب��M���������:W�ϖ����4�+�uW&������e}0���ו��� �!��ȼ����)PA޽;4�l����n짯�	,8�Q}����H���,>$�'f�ٵ�e�^˯ʹ��9���v�/���ml��9�r��}�����h��%��Xcbp��'輝��eN�ħƿ�9c�Ȋ;Gx�����W���5.M+S��<FΗ�͕�k!<�`�	Q!u��"��\#+��S�'���{+��"hac�'���Op�ե[�wc�}�![ǆ��J�>�&�����Op�ե[�wc�}�![t��ж`-�}.9P;��Op�ե[=�<r	Q�1r*:������٭>[ i朗-@IE�U����\u��\W��\�<�dQ*��P�+����&�D&���#�{�0;�}f�u�t��G��t��N��|�z��x���� �H|l"�n�)��W�sb�I�p\�WB.�?�����1����=��[,OV*�؂9� 4
���p,يg\#%%m�P�ŖmJHn��z�|=8�E<�l#�'�s��P{���.M^�% ��'��h�'���Xw�8����g�w�K-QS�)37J*u�,�JL���̀]�Bq,�7䔱+��TD��ό���.ӥq$�&GS�ГM��]�!��	Ǹ�y85��^�	 �wa(􆿳� w�6p�d�H9M\��e���S����g"�،j�����"��0��t����34�E����T��2$9]��ҋX����@�ڗe'x�< D]��7G#+�ǟ
��|�6|�+�� VU+I�z� dڃ�!�#��1G��LI�c�=��y�4�\���K�Q�]�(��X�7P��T��]�!���1����m��#l�p3�"�	[�*B�ﻋ-�����S8�����@!��P�h��]XT�g��U-�e5��e6²�/s�Ҥ�z��AqL�*�ﻋ-���C�M��N��SX1?�sE���ʹw�f6Sx�lޞ�ό���.���K�Qq�a>�WD���� ��'���Xwa'�<� \l�*(��'��Z���T�]�!���1����m�/s�Ҥ霁�q�0�/Őﻋ-���C�M��N��SX1?�sE�}��"�F2Sx�lޞ�ό���.���K�Qq�a>�W�0����'���Xwa'�<� \l�*(��'�"t�\˖��]�!���1����m���م*y=rJ���i3�ﻋ-��ȳ�Ǿ����n���4�$8�r��|0H#)�����R��#��� �:�����q9By�D$^�ggP��0��s�
��?wP� R��*z��y�+��W����@_Ϳ2�t%>^��7�ܥ��2��C��7�)�}�����T��.��W�������4:ˬ����Hx����ќ�
e���4述B���]zo}'�o�ee��&�dfl0���#�����Ź��������U-n�6j�+Q��΋|���.+ �I57���y�e� e8�~��(-��xsF�o��ǵ�ڊ�X3U�J��K}�n���?��}?�=\e��W��4�p(q�;�$�f�RҶ�ދ����!�]f��jI^�E�4i� e8�~��G$��"�֧z���>��RN#c�&ەF9#�[��ܶ������;vLď�C����h�MCTlS�ql�*(��'Ħ���aT������ e8�~����gľ�W���dx�b�W(��	!nR�K��AR%jg�Em���"B�䟷3��᧋�9ܧ!K��\4�.��jl���&�ى3ӿ,*�L��oI�] e8�~�� ��!~�2O�R�<�Uh�*�bh���d��f�`��X~�.H��@�H+_��͙�W��o?�`0��	yq�a>�W�7��� e8�~��<����B��B�BtQ���>Ft|�J �[�/����o��	���^�2}�0x����-Or�`�B�I&����,���s��r�m�V�����b�� e8�~���5��St4!=�)-�M���V�Yct(�P:��^��g��t�[9x%UOTmc���XYo�s�#��=�m�w�}��"�F2j2 |pD� e8�~��f��Ԡ8�tF���)e���n�`�v81⸟��0���x���"� (00�K;C�d*@��t�{�h�����#M;s5&��� Y�W@Җxh�Qf�h3Z6&�<�
e���4述B���]zo}'�o�ee��&�dfl0���#�����Ź��������U-n�6j�+�D���<\���~��Rʳ��y�e� e8�~��(-��xsF�o��ǵ�ڊ�X3U�J��K}�n���?��}?�=\e��W��4�p(q�;�$�f�RҶ�	����ܾ��.I"�т�L_f����@$˺/t��꫕qŧo��K�O�.
t�(XPrx�<�+��M���g$j�SX��{��ٴ��{�G��ͫ������:[ۚܖ��`�q�a>�W<�m=H!�7A<�SNp>�K���y�MON|�>�)5�(���{�eV���C�T��,�v:a����%L}pa��؊�"�D���al���:S=�]KW����@_Ϳ2�t%>^�߬Ҳш��?J	q솄|b!��u��Gɰ���:�#��:��L5ӥ���-���f����Oo;���6��B �ˇ
��lC��ۺ_~�M���g$j�SX��{��ٴ��{�G��ͫ������:[ۚܖ��`�q�a>�W�3�G���JA<�SNp>�K���y�MON|�>�)5�(���{�eV���C�T��,�v:a������!�=��؊�"�D���al���:S=�]KW����@_Ϳ2�t%>^�߬Ҳш��?�XQf�%~b!��u��Gɰ���:�#��:��L5ӥ���-���f����Oo;���6��B;���
ylC��ۺ_~�M���g$j�SX��{��ٴ��{�G��ͫ������:[ۚܖ��`��1Dg�Ŭ� �5�h�}�Cz���C�ҊQ �F��6%j_�z9�GKP�2�����Vcv�iL�D�"�
����Z�q�PO4�:_b�b2�����Vc2�����VcAQ@;�(V��6����|{��@�Pd	��0���3�R?�6��'�|,kW�A��ˮ��V�rsSRą���=]x�MԿǁ��2݆�?��xX0A./���d}��[�ƭM�]U��u݀�4h�t״$(�>g�qE�$ox�"��z�R ���ѡ�'	�?��[r(þAC#/<���qt�==�SD���Ju�Y��Ox9�t19@���.^Z�6^��<�b�؉͕$�;�N�C��_�~��xS�B7��A�hp�F�w��.�xI��v�5ܗus��t#��J��_�=�kM4v/��M��z-1�J�o�a�y����O�(f���5�r*Iީ�KY�`*y��	+D�}�w�k���9��:mh�a��v�cZ�Rh�|��w�Xb<�����a��xmlq�t��e�3DYB�*�+��.}��i7N�_��ϮD�R+d�8Dѕ	n�6��9�ȯ�ta;(XPrx��1�X�C�	�GݔO#�Z/��v
���M�wScpʎ/S�����k���9߅{ �����}��a�Gw�Xb<�����a��xm�%�緞�$r�t�}iV��	��y�'|:y#&�o}p�����:� �yD2�:{;�_��^��oF�:]�#�c+�g�0�u�1�G
�S�x?>�jޗ�	x H��em��գ��J,�/������>:&��~�K�x{^4��*m�S8�Lj�B�B���)����CF��f��x���Wh�x#�L_�(D{ͬ�y�4��������0+CZ�{9��K)>�=�������ʹw�f6bC4QC�ܯh�yy� �ˇ
��bC4QC��(�PF}�}��"�F2bC4QC�ܩ�`9߭�e���im�|���鉱�v\w�äa>*<UB3q�a>�W�d�ɏj�-M�O��~��ZD���A���Խc��J����WFIa�v��JaJ�1��� ��U�nFq�a>�W�+1,yՋ볺DLp�&�G��"O1����VPY���a	!33!�]f��js��pUo��;s5&��� �U��೧z׏�����M��|���5�ϼ�L��ߵ����h�1m<:E�pŤ'�]�a%��w
]�f���JD\zRc}w�M��1�t/ �ˇ
��۪	�}a�iQ��ׇ6�N�{��g{��Q3@�
�10�0�!�]f��jѝ|�+��X��WG ���H����宖�r 7
�8�
.���
�x(�i��/Rg�`�CB!�]f��jƜŏґp�H���ޓ���Y'"��V�Q��y���$}��"�F2{�R�$�V�q�a>�W{>����~:4�04�jf�,�(!��糳�huI�����;s5&��� ���Pf���x{^4��*m�S8�Lj��]�J��V����CF��	�Z�Y�h�x#�L_�h�:��p������"oS�E�� j����}#%�g8
����xQ�n
V~$q�a>�WȐ�-���
�2�z��v5���5ߧE4��Fi��|�),����2�����Vc2�����Vc2�����Vcv�iL�D��hK\K��h����V�ѕ���/����`9�GKP�2�����Vc2�����Vc2�����Vc�����=T��8��)��*��9�^�x�l��15�r*Iީ�l����h���X ���١9�G�O����	�B���y��z�U��&�Kp&Zc��g}Ю�0��%��	��@����!�;�Ӣ����a����C�|d����42�7g��zQ��X[MnQմ�u.'%vaA�E\���'�ZX^�O��N^�-�n�Lߩ���j��g�'���$k����#nn?lÝze�Nz4�\_G($�yܛ%��6�NHMI�!a$��OI�;�Жl:�������S,]G��wi���@�}z�vE��HT�����lf�%�B�>�9l\}=�ɕ�s�W�m/4@�s Oag���e��<6C¦��_�j?�N3�J�����5��gO�q�����f-#K�v]|nkظ�����or�}�!�5����04m��hF\�肬��2a�{:��so������d���aς"���@m����O��/D�_8\/Hi����s��.H'�t<9�	���K���9� g*"o�	t�F���U�K���K3��S#�F�K͕[y�;�Ӣ����L��1�gi�q���U��~�SA̃�����Z鎬����=���ޒC>?��@��mH_u.����I��w��,�\-�(��k�ND}K,��TD���rs�i��s�٭��[Ø�;�x\�HP@�a�b]�iz�y�Gs/�y;���\P+�}|��XH�����,>$K��(�+[�z)D�����pzl��a�d�l�gPk�c�z5�I�rs�i��s�٭��[Ø�;�x��`y���pzl��a�0�͏����c�z5�I�rs�i��s�٭��[Ø�;�x��`y���pzl��a�_����6Ƭ(Zy�뽑�,H@�Js�I��?t��yg����qu ��5K��~ҏ��Z��yt
cf�Q�-T�����Ps_*�GqW�w��fDB�	Kl�/�{u�_�%��ݞ�;a"U�T�/_��_��#g�k��CY� N��᧱f��:e"8���PyV��	��y'�0�U������;bЂ{z�0 �X��uU�v`,9�H�W��7s|�֣�w;��I��^���\�}��<P{���%���?����[�ˏ�����Z���삕�ռ:�4� ���?�Z�(v'�?���4��>.g��/�ciJ�y��ɩ��-�7���c�)�~>��hٔ9�ð��T�K:+>]�Dx���O�5ⰳ�-M�O��~Ӿ9�d�L�LT�;o����n�Ƶ�,0=]^	�&�2�T6���F3���%Ff"�	-7���RA�d><��F�^^d�3�-��&?z�	h�Qf��lա?mt}q^J=����x�ԉ�>B�R���>_:���!�#�<�  �ҋ�;#P�j2E�?�5ߧE4��c�}���Fo|k�Lbx(�i��/RŻ�&ǥ��4����m1�H���W�w��fD��<P{��Z�|��\�#�uf�8��m���`�֪���"�?�d���&��d��L_�G��U(%���x]�BF��������D�$0䅀��r�-~�$�1M�8���/��+!�|���l����4�n���xǊ�r"�ꉤ
�),`�LX��WG ��"Ҷ�ٔ��l�^9|�F�=�<�^�"L?����+�r5;%3���5(y��q9+t�}#k�˟ܒ�o|k�Lb��ܐ�}��JdT1�V��	��yQ��x�>'<!P�:-醁c�����*_ #��P��Ӛm��{%檛��BJN��{~�@�i7N�_�ߑʰӔܻ�J���Z���,�j8�p��<���
f���P'��}���^���\�}g?	��o�׵���\"��6,{�0h�5e��y���t�T���"�a�I�q�����1Dg�Ŭ<���Hn
V~$����)�V@&� ��LI/��\]��a-6�Da�o�eC
�Fk_���F<���Hn
V~$��S	���`g��%��v���q�)]Q�x��r_��m�,�j8�p�V8��R'�U�4M:1ǃ|	s��#P�j2E�?�5ߧE4��c�}���Fo|k�Lbx(�i��/RŻ�&ǥ��4����m1�H���W�w��fD����r�- b��)j���,�j8�p�0��ܗ�
f���P'#�
_�jE^���\�}g?	��o�׵���\"��6,{�0h�5e��y���t�T���"�a�I�q�����1Dg�Ŭ<���Hn
V~$����)�V@&� ��LI/��\]��a-6�Da�o�eC
�Fk_���F<���Hn
V~$��S	�B��w%��v���q�)]Q�x�p�NX9V�3���5(y�<���Hn
V~$��S	�B��w��,��>�,y�Xi�A4^���EqJ�1��씑�:��KY׏�����Mrw�&�z<aSm�6��`߸��S�Ȍ�>>Y�k9;��|B������0��ܗ�
�E�i�m}66j�"Hs���S,(�<�/�#[��$�M��j��p�Ե%����r�-���~�ul����4ۨ႑9����O�sL~΄gO�3f��*��������[�/O!坭�悬��2a�{:��so�9#T'��nҍ	g�y���5��gO�q�����f-|�bxKҲ��r�D� �m�'4�a��䒟JƓ����i�!54�:esĘ>��F^aQ��O�O�d��e��C}��W0i��^#j#ổ���.D7�G�Ai���KIF���%�u'���Xw�j�7���˷���T�\ �͘�f��p�b�z'hۉ)��R��삸1Dg�Ŭ��{l�f|�ό���.Ә�ʤ+�+t������1'���Xw�����U�fY��Up��m� �˟Z鎬����=���ޒC>�W�~'D�i�l�u��]�!���\B��VPg�2���� b�@IE�U����\u��\W��\�<�dQth	 ��T���&���#�{�0;�}Q�; ��
*�+�i�0� V��I��A>��d�٣��c�A�L'������"X��[Y��kB�h=Q�Taz@mA�^,�V5+��:�g�ծ,��[Ø�;�x��˚����Z��LA�w1�;��܇I�t׋Q��Q�E�%�i��;��|B�M%>Y%��]}ҭ�gjZ��s_4��>.g��/�ciJ�y��ɩ��-�7���c�)�~>��hٔ9�ð��T�K:+>�~vBc$׃]��+5u-M�O��~Ӿ9�d�L�� l��'t(�aN��/X��WG ���e>�aq�cY���R�Ĥ��	�_]���n�#�ܮ�E���7t��"L?���/V�/��Y���j��ܒ�o�r:���ní&���.�Ȓ�p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb��ܐ�}��JdT1�V��	��yh>Q`PQ�{9���LA�w1�;�/����G��C0k���%�i��;��|B�M%>Y%��]}ҭ�gjZ��s_4��>.g��/�ciJ�y��ɩ��-�7���c�)�~>��hٔ9�ð��T�K:+>�~vBc$׃]��+5u-M�O��~Ӿ9�d�L�� l��'t(�aN��/X��WG ���e>�aq>ν3�`����#�4� �4�D7�@�B�xȀ��D�[b%Ɨ�����a�c��9"�0��1Cc׶
�b�]��xȀ��D׏�����Mp�-a�D͢q��`�L�5ߧE4������!2�͞nOY��G�Ȧj��}jj+^��z{�0s��O�h�	?�d���&�L:v�
XJZ��S$v�0�x ��0��1CcכeSd�̣�_2��VU(��z�j`0��a�S����cܺ���T�Ѿ��/@�&����`w�:�%��R��cՇ���J�NId�p ~��Z2��R\B/[͋Ip��}K��kظ�����or�}�!�5��Z�T1ۂ�r���x�d��䖯��l����4$��p`Ԡ�U��%S�;���Ų���(i.ْl��]�B����&�b��_�G��G�^ֻ����XP��ȟ^+r��C�'$�7g�@�;ۂ��IÙ=�H9�|!�4����?`���HH
�2y����#��v�~������]�!��	Ǹ�y85���s#%��"X��[����fbK7͍��|��W&":�AuFT���č�Y���S�)37J*u����8d���u�"�|��].��'���Xw�X�����Z�oO�q����{l�f|�ό���.��W�D�b�v�~������]�!��j���f{ �$���{l�f|�ό���.����`4�E%v�~������]�!��E��}��n��9�n��(�
t�������2�b]�iz�R��G0�6�������-�@��X��H��*֪r��C@�19&xc闑^�$��Xo�`��]�E$��*��b�JHn��z�N��xo6�Q�J�V���1��I�:����Mׇ5����`K�����svfY������^ֻ����XP���	�$��ɍjώ�au�0�cܤy䓓ʉ�8�!�I�<�[[B�����'���Xwd�n]N���k��i�qs����R�wX��\o�LCd�ĸ>@��H�`�-�IBo�A;h�F$�Μ��VK��!�O���E���T�	\����]x�l�I��R�ﻋ-���>��l%i�-b!��u�>���6���[B�����'���Xwd�n]N�\���dC��@����	a(􆿳�"Ǝ��_���.JL |�7J����� �!�( ��@��7� �91o6{DPf_����g��)G�J�cbp��'@
9��y�	��F|.!h�67���	� 1��=ە��ز�FFh��Wǖg3ȓ8���/����h�99φ��<�6�����b�s������cp6Dq��;���EWr<�_�/_G��'n�^0o**�ХM
�NAJkD�̆h�67�G<��N:h���8-|�D�H������@�0�.�����/d��-����G����?�6" �f:^օ?D^���zg��p��+p����,��nF���<�W�.�P�	��
�Q�}�����!�`�(i3)'�{u@������h�Ш怛�6U�.P	HȆ�?�Q�9^�����hg�d�H�RtV�^!�`�(i3r���[��X�Ղ����<���H1tSjv�!�`�(i3����l��ܯ�.ȚJ����oJ���9�i	A��Z���Ӗ��x�?�+��d��MT�scX{�X!,!�`�(i3G����?�6" �f:ҭuF,!�`�(i3�ʥP��e:�K�PP����.��N�!�`�(i3!�`�(i3��jVѭ@!�`�(i3!�`�(i3԰_���{»�A\���6" �f:����M�!�`�(i3
�:qEp�;�P�t�5!�`�(i3!�`�(i3ܩ�9�d$�X�⺘EBv�@W&�g9���.:��Q?M8�f2!�`�(i3!�`�(i3����fE_7��C��k����FrTA^R�v0 ��??����}Dq�f�!�`�(i3�zg��p���of\m0��#��J^��҉�O��m��J!�`�(i3!�`�(i3�u��A�0���򴶽!!�`�(i3��w�w:�!�`�(i3!�`�(i3� ��D�	��!�<�����ć�8���/��z�V�҆�7�j�e��11�g��U-�e��,H/��!�`�(i3ʐ���~�T��0�����͖n�\�b��\����`��!�`�(i3$f��_Ub�F�S�1 �
�:qEp�;�P�t�5!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�׹��L<C%`��L�b�Q����,�4�Ŝ҇���e�(B��