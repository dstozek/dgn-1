��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t����j�X�8�����$4L�������}g7l�� *��I������,0�z8O� ��t'�O��!y}_���C���cC&��BB�m����_�2rI~�K0�HR3=�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K�ų��/���_�^�r6}F���XTcFǲ�r�t[e7l^�Eu�n�=�"X�崺%����ή�6V$4���,-O��0:��(5���]������[��/1��-�F�	G�ಥ�}��၈��`�s�smyo��9��5�ܧ6�(1E��
�����ɸ�Bo�Uޣ���]�9��2�@�� �,���S�8�I6�qB�j����iҕ>�>SEV�����[�t(D�0��g�@��\��6q*�P��sz�֛����w�W�Ԇ�9�ޑ�L�)�܌��F��6D%�4�v�������h(`SR'k����Te#���VtB��.�����(S��k`5���7���j<ҝ��R��,�vzd���Mx4���x~`� dȜ�^q2h�ڥS4�}eױH�;��k�/�꠬g��h����Sǘ��� ��>[I���d��{�Jl�Z�PG�gx��3)C}��;1q:���?"�&����\���	XӈjB���IU{Q=W�]3�ǧoj'í�S��z�}���HJ����5؎�T�(�#�6���h�����of��C��l�@	�nc���Rp�YX���H�k�e�w΂�9~}�V�
���W���T�MNU������V?`Tӓ�>gA$��4ѣ �ؓ�=6��}ئ�X&]�����Ӹ�H���E�^�0�x�t-��ϻ_4YwA��r�l+^H���v���ƺJ�ٞ��x����e�A�;����Bk��2�,���y�U�"������)��\3�*�H(�Bd:^L�:��g$b�̦� |)_3��3�@D��d��Ǉ�Z�}v��ى�\I��g�0��_�o%�����L��TO	w�ǆ p�Ai�u�1mv\�[ak0y��/�S�a�1�����@��F0��|>�a�,���^'Um��7�ΫjK��C0u��{������+�X}�cE������܆N���l���HZ��>�7Jjb`�h܅
��0'p�P6~&7z�t���+�m�(R//|�X�5��*ꊞʮ;����kM��WIkH�ӯ;�@(�}�t��m'.�����0E�ڔԱ`��|M΄��Z �r�M7tL>z��Ux>Fs�<a�J�WЄW����,K�H����ނ�6t�+(�1�uf�G�5���zr�xЏ��|�#��c�Mp����Bv�-��`�g�t	�W �{}��(q 	�����g�����&�a�T�=�q<.BLN3�
Cj�fU�A8ܓM�5q~��nH8���L�òfHS���&)�"�<*�Y��nZ�)~�%�����ʽ{�w� `j������>�DSA�c����H��׶�faΉ{�M���CQp
s2��z�؜d=a�3���C��#��F�5P�I2]]�������������;�z�h�D���+��8�[#�le��2TfC��(n��L��=@Vݺ�t�DЮ6��c��J]y��|.��Lle�5t׶��-�M�a�Ҹ���"G��(�M�����(ĉ�jZ� P_࠶��4�a�����!��� ��Ո7(p%��0hƵ�S��29@��������>��h����V�1z�f�{\��i���,K�N`���Xsw�M����·
���
��O�z>g�Tb8<���y�F����\��T��	�h�UN��.�M$�^��O����<	>��PN�;X��H`����v��q�._1��ޠI���y�^c�4��}Ժcx��Ni�y� Jf߳�8y�y+MH><g �H4\/�7O��k)���u�I]Ai\DYg�x��,����I������$��b��a w�$��lk�pr�F�D0����>c6R�1�_���󠖩*��5
��Q�t��ɨŹJ=.��h��� 2[�KfbM��ȓL�S����TS��})z/�(u�H���g��VD+a�-����F���\� �#~QHP{��[�H�%�P޸(���d�px�7�Q��!���,�ȓ=�藧Â(�c���l<Jÿ��o^���: �T�@Z"#�~���K)eZ(�S8%�S�P��֔t@�1��@�\�nZ������F�i�	D�ͦ	q�c2ApG�p"6%����i�@i�š#yyY���O*3��Z;�5#: <�]�2{+����Mb�mtY����Gw��. ����݂�K��6�V�������%Ҭ�}�/���h����ZK���0����6�[��~��F�\��P��B[H��QX��X_���f�m����h��B�p�5-ݔ�m��Z�׹��g��ކs$�NѪ�ʅ�0>d�Ҳ��?|y��t�Uwlj� J۸�м�i���V�7E7��a�F����*�B���h;A$;�K�"�ҙ�"�&P+ٹ���b�Fx��H�w�����D1Ђ�C|T;ڊ;�M;�	�8�>���a�� �i���>���<��
�{YՖ�M�P�r�sK�.M��_,h����$�_YiΛjki?ԮI�1��B���=��<����U&+�����]�x�F��5�Q��d^�ȿu�'+K�7 B��Vx��F��@Hn�P&c��zK�V��Z}'8��0�n� �<R��h"���i.@]b�I�;�wbn���1�0o�Ϟd� �r�o���<�XqeY�r��?/�l����^��O���HC��ٮ$½�e�r��ϣ�X�x�i�L�5@w��[F�T���TS��rp�JuNd/��^��S�]�c����t�&ϣy5�!,�Q݇���z~3���{�u�K��(w��8J�|@�,�\1J%�e��Ņ"U|묂�;�����_pт):ś�6b�.�ɶh�⠮K��<JÀt{,�ރ56�������+�f�Ƭ��� ��&��v�U�f]��O�t�5V�t�����W[�'T��I�9�i"��4Z��N��X�̔�M+��R�~� ��|���ʇ���UF��5�S;󕔟�b�I�ˣ��x`>���C��u���P�s���©�z���i���6.�ďJ3���y�Kŀݝ6cr#�=�h2�{�jar�ч�QY�ES���3cP�|b1�[]�$R�����ps'��	�
�8�m�3L]S4��w��51�\0�2M�\`ŖA={=��#��*�� 6(}W,T�%c���[�R�e�,3��Z��� �ƣbQ9��᫣�S��