��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t����j�X�8�����$4L�������}g7l�� *��I������,0�z8O� ��t'�O��!y}_���C���cC&��BB�m����_�2rI~�K0�HR3=�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K+Ke%G���N�;5LR��>7���F�dR�;�#a�=�?�c�=m#����?�5�^���f+ns�����
��%p�2�P��}��'!*b�6�H��V%wX��oܲ���|9�F >��T��ކ)f�`q��'����O:��u�-����Z:�eN�[��d����.}[�S�H����o8Z�e�� a�]�;���^��W(W�9ɏo����CU��k���^!�5R@�zU>�&�i�C�(�p/u���&��NI�5�ض���G�q8���I^��J�Ll�#/�W��	�\��ks�\�w�*��:�3�U��W8 ����T��(���r@l4�v� jp1�I�'W��I��bo��K'��ʸ��\1?���d{{��,�@T��Zj��
�n/�c/Ɖ�Eȳy	���,a,?��M���1DW}��7�����!�9��E$�=ڝ�J�1$���ء���R�.`�d�#h�S�vĘ�0vtMw�������`,Ţ�$�Q�
�Ϯ���K*�Ȕ��X(�!P �#�˴0�����a����=���R�y�Hsu�p���e�:7�v̜�Pd�txv⏵����A��t�l
Yd:)�K�������U��u�5�(�9�;��]�pK��:R��~	����~��.CZG��G�.��,-������ʆ8�K��f�̍�`�@Qf��@mH�sک�"�C������v�ܢ�M0�;�3�������d���L1��=��z"?���0����,�gQ��<jR*Ǝ~C�a���oA[7���wS�M7����C��:�C�N�E#!�"w�z��1a�!u�����ݦ�Yc���-��g�E<U�P$��"��g���0"K*�V]�S�)S��b{j���du�)>�:��-U���[�tx5&=C�^;��k�� �]�7;%� �.�hj��������ю��p�J�ԩ���!�{��u*)u�g�WKg&�ڦ��Ih���3E£�$#�w����~dIY?)�|KKD�y��� ��=z?=7���7��Oe�7�z`c��j�Z�JFN��[-xQ��ͺ�Dp
}<j<���"5�RdLNթ��Y�J�C����C,�׊:�LArR�{������W�+������RnI�x���s�����W��c]��+�Ʌ�����8�O'��Z]����ݝS,��� n��� >�h��U����\���	�[�\I������ٍSc��L7�����+�G����?��w��.�����~�7��nBB��
�sL�Wm�чp�)Ǩ0^���%���z<�'��K���F�
T�@Gx�)Y�����O�$��b�wU_�$�Ũ����_kL�+9Jػ���	'tЈb��zs��jVq�f��E\��Z���9����m����O]'���˻"�UO�R�GY���ֵ绝N#�D�� ��.���+@�C/��F��V��V�R�����T���1�R� St���̄y�6:�Vg���Ӣ:d[�tR��x�Cs�1z��΢y)��L�PH��L.������:��U]ƹdx��
�(�/8=\E��Y�o�>G{�ۭ8�M(��;�Vxn)�%����f/0�0������"1U��8�)�1yw�9�q��$�%q��}m��y3�?�ቇY)SՎ�1��s�,�5��n/���|g�����]/��2L���_�lK��e�q,3��Q"�68U\y׌7�e��G`8��6h�|��@#��XhG��)3��Rxz?�����fq�9��9��Z�+ir,�s���-}M�F�@m���ϝ�E�"�=!}/,��j ��<%I `{-�Q	`>(�=vǁ�d�H�br�0.�^{W�Ou����8� ����[�B�u�� <$R�o�\Yjw��������@�P>���5�f:��3D�Ղd�a�i��"MK���e3���_5�ʝ^���^L��N�a�z�Lq%�=�0wQZjk�ŐVG��4�۴�$��C�/��� �ل�ax2Ntj���|4�2-�����r��orU�N�8��l��l���+��OǴ��b5�:�驶�>��*U��G��R,l�ɷy�is����X���h�˫s�Q�͔TOK���jR�����$*�9�I�#f#��h�R����ci�?�]�d�\[���t��)pRΜ-Fp�.C����Z*��P�G�C9K�m��r��r�̋M���� �}�p�}:��Q�E͖��l�<�/d�8��جl�ߢ�[jfemY��]��T�&�k\�@���gm[E��_��ݰ�X��_���C۽���-�	�������|�T�E���0�e�q�Z�4ԉ�����+�ܶ쓞u8Rb0�SLv���Q��º�Ѽ�Y�C��gԷ�����j{��m7˯�82-��XZ�͚�.��G���k}�gP�1J�mߔ��j�>Q&Ә[bN�Mc�����[�֮�/�-4�v7���_c�?E������QJ붺��J����}�ڪ��yP6��JWWBl��1�*`����O!����0(�	G {���������2�*�T�<[^��1LB�?�Z��h>)i{�k�BM�4��ODz=������צ���pcřVd`!�����1*^~`���E����P2+*���tr�7R���tǒkۋI�|+���-Ώ-F�s�,D������ړ�^צ�����%V`�?�lU��P&���S6�t�G�O���Va��w�Sd�OʼO�����|ݩ����H���d u-�;}+���Y�*���Z�.+��N��D�)�����Ʊ��{`�A���f5���u���:��u7Y�Q�yv.�9\�_��LHˠ[�/�w��B�G��������f��#V�0���;l��Z�'4�:�6G�g��lЛ-�.�s��6�<Z�e��-R�yO5UV�EF��7��td¾�U����'�����34����hC㒆��Z�K��)��Sl+8s�m;�&-�5��k@���rs��8H"�c�=`��4�c�yLP�� +M��=�'㌨"��'�"%nx���',��@����ʁ�o*[�%��WS7�c��m')��L�$�2��U~������`Q��5Ͽ��
M������E�	�i @֕�[bdiP��"��`&VN�O
���-��J<���;
�[2oߴd�(@�O`M���~�Jk�uì�6����S�����Xg�P��4�4Ƣ�N8�6L\] �I��l��qbu T��Y�#]�#���m
�m���X���c#��҆X1X�A����_k3��-$�}rU�!���ԉ'�9����:$���NSX}
�$���Z������F#����[4����B#{m
��{��Ɗ�{�*�%~����v��URĔ���Re�ͧg��/S��-�S��N~�M�~�� ����F�D���	o���@/���,��W&��
��
�:>�鏒��8��nM�Z���f�<k�j�G����x�y#R�n=UH�WM�"���54p�T#R>�^�����`��N�c>O��=��m
!����7��⨂���=hy��|�W���_��ĈУ�?���٭e[q��&�z�:�R(�U*̄v����qiJ(y�Ɇ��c@�MN���G�ؒ^�]4ʨ�ƈ/2k�#�	��Uh�p-'���uI;y& 𐱇b����}� *l��@u�Ĩ�k"�|�J���_u�ⷱ��VM"�GԄ��TTY�.kV[�1����`�_L�;<��ל�͟"
���Ц�/	Y�*�Z��.�� l�=
��%�{���U���;~+��]ۍ-�N���iU���زH[�i	���kI-�$�$7�m��2B����$Z�!�T���13�a�2�]j�Q��@t�2�*�p5�_��2Q���\��eJ�9ŭhL�]��xW�Qձ��%a��A���e�૯36S�����O�&v�A;��eI��SkV�"}�7![?�e����0�������Љ�� q��Q
Z���4�{��u��;�h!ڽ��̜.�D��q��u���c8 3,R4�Mb�G����]qv߱��!�O�#VPl�p���$;��j.͝�c���iKN:�IROt�{��t|�����b}-Շ�mM~1��-K+��<o?��j��*��DG�ήEZ$66�9�
���=>rUq�1
�����Yk,��#���qb�xȦ�Ք�@|DQ&}յ��DmZ ֖@U}K�3�n��K>
�م�"1Q��������F��IJZ\�/��1�yk���U��Z/������BF����'���Q�����@ﳟ\<��䟢��k5l
K�ӊ���w�Q#75��h��n_F��mH�:�?���z����s��a��sE�0�'��K��ȕ���;n'�%=��B�w���qU8��j22�2�'��U�p�z�|�~-�NE�:-��^�(O����������l2X���:J��/%�x��w�L����9� U0�Yă'�&�#��{�U*H�0eɂ��0L�ɹ�N'3�n�i��*�ԉ�O
.��+_J���w�PR���^�`!��gag����WXڔD:	�R��5n��bq�5��\@�;��gf���Ǔ�������&:�B�b	%�v�
wgQ�A�@Y�t��3��]n��.6�Q�����g<�!����10`��ٍc�m��š]��k��'��t%|H�zG ����Ӣ��Aj��������R� ����A�Fl�{�a�)[Q�㌿�%��?28���/�Ǹ���s&"��s G���E��+���.���W�OvCq:�؍��@�<dk*e!�Q����/�������Aե4TNnF�)�
���i��l՝�婆=�rq)(��]��,�q@ �L~JC�'r��XO���K��zz;}}f�SK�f��!�ܤz��Z��c9�