--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arbitrator is 
        port (
              -- inputs:
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                 signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                 signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer : OUT STD_LOGIC
              );
end entity Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arbitrator;


architecture europa of Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arbitrator is
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_allgrants :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_allow_new_arb_cycle :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_continuerequest :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_counter_enable :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_beginbursttransfer_internal :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_begins_xfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_firsttransfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_grant_vector :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_read_cycle :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_write_cycle :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_master_qreq_vector :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_non_bursting_master_requests :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reg_firsttransfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable2 :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_unreg_firsttransfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_read :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_write :  STD_LOGIC;
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa :  STD_LOGIC;
                signal internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal shifted_address_to_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer;
    end if;

  end process;

  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data);
  --assign Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa = Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata;
  internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 22) & std_logic_vector'("0000000000000000000000")) = std_logic_vector'("100000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa = Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter set values, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_set_values <= std_logic_vector'("001");
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_non_bursting_master_requests mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_non_bursting_master_requests <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_bursting_master_saved_grant mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_bursting_master_saved_grant <= std_logic'('0');
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter_next_value assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_allgrants all slave grants, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_allgrants <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_grant_vector;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer <= NOT ((Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_read OR Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_write));
  --end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer AND (((NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter arbitration counter enable, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_allgrants)) OR ((end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_non_bursting_master_requests));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_counter_enable) = '1' then 
        Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_master_qreq_vector AND end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data)) OR ((end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_non_bursting_master_requests)))) = '1' then 
        Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable <= or_reduce(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_data arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable2 <= or_reduce(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arb_share_counter_next_value);
  --cpu/data_master Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_data arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_continuerequest at least one master continues requesting, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND NOT ((((cpu_data_master_read AND (NOT cpu_data_master_waitrequest))) OR (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write))));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data;
  --cpu/data_master saved-grant Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_data, which is an e_assign
  cpu_data_master_saved_grant_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data;
  --allow new arb cycle for Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_data, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_master_qreq_vector <= std_logic'('1');
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n <= reset_n;
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_firsttransfer first transaction, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_firsttransfer <= A_WE_StdLogic((std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_begins_xfer) = '1'), Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_unreg_firsttransfer, Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reg_firsttransfer);
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_unreg_firsttransfer first transaction, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_unreg_firsttransfer <= NOT ((Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_slavearbiterlockenable AND Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_any_continuerequest));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_begins_xfer) = '1' then 
        Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reg_firsttransfer <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_beginbursttransfer_internal <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_begins_xfer;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read assignment, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND cpu_data_master_read;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write assignment, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND cpu_data_master_write;
  shifted_address_to_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address <= A_EXT (A_SRL(shifted_address_to_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 20);
  --d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer;
    end if;

  end process;

  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_read in a cycle, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_read <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_read_cycle AND internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_read_cycle assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_read_cycle <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_read_cycle;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_write in a cycle, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waits_for_write <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_write_cycle AND internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_write_cycle assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_write_cycle <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_in_a_write_cycle;
  wait_for_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_counter <= std_logic'('0');
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable byte enable port mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa <= internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa;
  --vhdl renameroo for output signals
  cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data;
  --vhdl renameroo for output signals
  cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data;
--synthesis translate_off
    --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_data enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arbitrator is 
        port (
              -- inputs:
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write : OUT STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                 signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                 signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer : OUT STD_LOGIC
              );
end entity Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arbitrator;


architecture europa of Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arbitrator is
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_allgrants :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_allow_new_arb_cycle :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_bursting_master_saved_grant :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_continuerequest :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_counter_enable :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_beginbursttransfer_internal :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_begins_xfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_firsttransfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_grant_vector :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_read_cycle :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_write_cycle :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_master_qreq_vector :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_non_bursting_master_requests :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_reg_firsttransfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable2 :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_unreg_firsttransfer :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_read :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_write :  STD_LOGIC;
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa :  STD_LOGIC;
                signal internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal shifted_address_to_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer;
    end if;

  end process;

  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control);
  --assign Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa = Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata;
  internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 2) & std_logic_vector'("00")) = std_logic_vector'("110100000011000111111000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa = Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter set values, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_set_values <= std_logic_vector'("001");
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_non_bursting_master_requests mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_non_bursting_master_requests <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_bursting_master_saved_grant mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_bursting_master_saved_grant <= std_logic'('0');
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter_next_value assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_allgrants all slave grants, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_allgrants <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_grant_vector;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer <= NOT ((Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_read OR Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_write));
  --end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer AND (((NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter arbitration counter enable, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_counter_enable <= ((end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_allgrants)) OR ((end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_non_bursting_master_requests));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_counter_enable) = '1' then 
        Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_master_qreq_vector AND end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control)) OR ((end_xfer_arb_share_counter_term_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_non_bursting_master_requests)))) = '1' then 
        Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable <= or_reduce(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_erase_control arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable2 <= or_reduce(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arb_share_counter_next_value);
  --cpu/data_master Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_erase_control arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_continuerequest at least one master continues requesting, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND NOT ((((cpu_data_master_read AND (NOT cpu_data_master_waitrequest))) OR (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write))));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control;
  --cpu/data_master saved-grant Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_erase_control, which is an e_assign
  cpu_data_master_saved_grant_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control;
  --allow new arb cycle for Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_erase_control, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_master_qreq_vector <= std_logic'('1');
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_firsttransfer first transaction, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_firsttransfer <= A_WE_StdLogic((std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_begins_xfer) = '1'), Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_unreg_firsttransfer, Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_reg_firsttransfer);
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_unreg_firsttransfer first transaction, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_unreg_firsttransfer <= NOT ((Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_slavearbiterlockenable AND Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_any_continuerequest));
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_begins_xfer) = '1' then 
        Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_reg_firsttransfer <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_beginbursttransfer_internal begin burst transfer, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_beginbursttransfer_internal <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_begins_xfer;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read assignment, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND cpu_data_master_read;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write assignment, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND cpu_data_master_write;
  shifted_address_to_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer;
    end if;

  end process;

  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_read in a cycle, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_read <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_read_cycle AND internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_read_cycle assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_read_cycle <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_read_cycle;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_write in a cycle, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waits_for_write <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_write_cycle AND internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa;
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_write_cycle assignment, which is an e_assign
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_write_cycle <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_in_a_write_cycle;
  wait_for_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_counter <= std_logic'('0');
  --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable byte enable port mux, which is an e_mux
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa <= internal_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa;
  --vhdl renameroo for output signals
  cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= internal_cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= internal_cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control;
  --vhdl renameroo for output signals
  cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control <= internal_cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control;
--synthesis translate_off
    --Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0/flash_erase_control enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity alpha_blending_avalon_background_sink_arbitrator is 
        port (
              -- inputs:
                 signal alpha_blending_avalon_background_sink_ready : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_source_endofpacket : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_source_startofpacket : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_source_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal alpha_blending_avalon_background_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal alpha_blending_avalon_background_sink_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal alpha_blending_avalon_background_sink_endofpacket : OUT STD_LOGIC;
                 signal alpha_blending_avalon_background_sink_ready_from_sa : OUT STD_LOGIC;
                 signal alpha_blending_avalon_background_sink_startofpacket : OUT STD_LOGIC;
                 signal alpha_blending_avalon_background_sink_valid : OUT STD_LOGIC
              );
end entity alpha_blending_avalon_background_sink_arbitrator;


architecture europa of alpha_blending_avalon_background_sink_arbitrator is

begin

  --mux alpha_blending_avalon_background_sink_data, which is an e_mux
  alpha_blending_avalon_background_sink_data <= pixel_buffer_avalon_pixel_buffer_source_data;
  --mux alpha_blending_avalon_background_sink_empty, which is an e_mux
  alpha_blending_avalon_background_sink_empty <= pixel_buffer_avalon_pixel_buffer_source_empty;
  --mux alpha_blending_avalon_background_sink_endofpacket, which is an e_mux
  alpha_blending_avalon_background_sink_endofpacket <= pixel_buffer_avalon_pixel_buffer_source_endofpacket;
  --assign alpha_blending_avalon_background_sink_ready_from_sa = alpha_blending_avalon_background_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  alpha_blending_avalon_background_sink_ready_from_sa <= alpha_blending_avalon_background_sink_ready;
  --mux alpha_blending_avalon_background_sink_startofpacket, which is an e_mux
  alpha_blending_avalon_background_sink_startofpacket <= pixel_buffer_avalon_pixel_buffer_source_startofpacket;
  --mux alpha_blending_avalon_background_sink_valid, which is an e_mux
  alpha_blending_avalon_background_sink_valid <= pixel_buffer_avalon_pixel_buffer_source_valid;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity alpha_blending_avalon_foreground_sink_arbitrator is 
        port (
              -- inputs:
                 signal alpha_blending_avalon_foreground_sink_ready : IN STD_LOGIC;
                 signal character_buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                 signal character_buffer_avalon_char_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal character_buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                 signal character_buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                 signal character_buffer_avalon_char_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal alpha_blending_avalon_foreground_sink_data : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
                 signal alpha_blending_avalon_foreground_sink_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal alpha_blending_avalon_foreground_sink_endofpacket : OUT STD_LOGIC;
                 signal alpha_blending_avalon_foreground_sink_ready_from_sa : OUT STD_LOGIC;
                 signal alpha_blending_avalon_foreground_sink_reset : OUT STD_LOGIC;
                 signal alpha_blending_avalon_foreground_sink_startofpacket : OUT STD_LOGIC;
                 signal alpha_blending_avalon_foreground_sink_valid : OUT STD_LOGIC
              );
end entity alpha_blending_avalon_foreground_sink_arbitrator;


architecture europa of alpha_blending_avalon_foreground_sink_arbitrator is

begin

  --mux alpha_blending_avalon_foreground_sink_data, which is an e_mux
  alpha_blending_avalon_foreground_sink_data <= character_buffer_avalon_char_source_data;
  --mux alpha_blending_avalon_foreground_sink_empty, which is an e_mux
  alpha_blending_avalon_foreground_sink_empty <= character_buffer_avalon_char_source_empty;
  --mux alpha_blending_avalon_foreground_sink_endofpacket, which is an e_mux
  alpha_blending_avalon_foreground_sink_endofpacket <= character_buffer_avalon_char_source_endofpacket;
  --assign alpha_blending_avalon_foreground_sink_ready_from_sa = alpha_blending_avalon_foreground_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  alpha_blending_avalon_foreground_sink_ready_from_sa <= alpha_blending_avalon_foreground_sink_ready;
  --mux alpha_blending_avalon_foreground_sink_startofpacket, which is an e_mux
  alpha_blending_avalon_foreground_sink_startofpacket <= character_buffer_avalon_char_source_startofpacket;
  --mux alpha_blending_avalon_foreground_sink_valid, which is an e_mux
  alpha_blending_avalon_foreground_sink_valid <= character_buffer_avalon_char_source_valid;
  --~alpha_blending_avalon_foreground_sink_reset assignment, which is an e_assign
  alpha_blending_avalon_foreground_sink_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity alpha_blending_avalon_blended_source_arbitrator is 
        port (
              -- inputs:
                 signal alpha_blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal alpha_blending_avalon_blended_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal alpha_blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                 signal alpha_blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                 signal alpha_blending_avalon_blended_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal vga_avalon_vga_sink_ready_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal alpha_blending_avalon_blended_source_ready : OUT STD_LOGIC
              );
end entity alpha_blending_avalon_blended_source_arbitrator;


architecture europa of alpha_blending_avalon_blended_source_arbitrator is

begin

  --mux alpha_blending_avalon_blended_source_ready, which is an e_mux
  alpha_blending_avalon_blended_source_ready <= vga_avalon_vga_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity analyzer_input_left_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal analyzer_input_left_avalon_slave_readdata : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal analyzer_input_left_avalon_slave_read : OUT STD_LOGIC;
                 signal analyzer_input_left_avalon_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
                 signal analyzer_input_left_avalon_slave_reset_n : OUT STD_LOGIC;
                 signal cpu_data_master_granted_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                 signal d1_analyzer_input_left_avalon_slave_end_xfer : OUT STD_LOGIC
              );
end entity analyzer_input_left_avalon_slave_arbitrator;


architecture europa of analyzer_input_left_avalon_slave_arbitrator is
                signal analyzer_input_left_avalon_slave_allgrants :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal analyzer_input_left_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal analyzer_input_left_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal analyzer_input_left_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_begins_xfer :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_end_xfer :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_firsttransfer :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_grant_vector :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_in_a_read_cycle :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_in_a_write_cycle :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_master_qreq_vector :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_waits_for_read :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_waits_for_write :  STD_LOGIC;
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal shifted_address_to_analyzer_input_left_avalon_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_analyzer_input_left_avalon_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT analyzer_input_left_avalon_slave_end_xfer;
    end if;

  end process;

  analyzer_input_left_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_analyzer_input_left_avalon_slave);
  --assign analyzer_input_left_avalon_slave_readdata_from_sa = analyzer_input_left_avalon_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  analyzer_input_left_avalon_slave_readdata_from_sa <= analyzer_input_left_avalon_slave_readdata;
  internal_cpu_data_master_requests_analyzer_input_left_avalon_slave <= ((to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000110010000")))) AND ((cpu_data_master_read OR cpu_data_master_write)))) AND cpu_data_master_read;
  --analyzer_input_left_avalon_slave_arb_share_counter set values, which is an e_mux
  analyzer_input_left_avalon_slave_arb_share_set_values <= std_logic_vector'("001");
  --analyzer_input_left_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  analyzer_input_left_avalon_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_analyzer_input_left_avalon_slave;
  --analyzer_input_left_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  analyzer_input_left_avalon_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --analyzer_input_left_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  analyzer_input_left_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(analyzer_input_left_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (analyzer_input_left_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(analyzer_input_left_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (analyzer_input_left_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --analyzer_input_left_avalon_slave_allgrants all slave grants, which is an e_mux
  analyzer_input_left_avalon_slave_allgrants <= analyzer_input_left_avalon_slave_grant_vector;
  --analyzer_input_left_avalon_slave_end_xfer assignment, which is an e_assign
  analyzer_input_left_avalon_slave_end_xfer <= NOT ((analyzer_input_left_avalon_slave_waits_for_read OR analyzer_input_left_avalon_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_analyzer_input_left_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_analyzer_input_left_avalon_slave <= analyzer_input_left_avalon_slave_end_xfer AND (((NOT analyzer_input_left_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --analyzer_input_left_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  analyzer_input_left_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_analyzer_input_left_avalon_slave AND analyzer_input_left_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_analyzer_input_left_avalon_slave AND NOT analyzer_input_left_avalon_slave_non_bursting_master_requests));
  --analyzer_input_left_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      analyzer_input_left_avalon_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(analyzer_input_left_avalon_slave_arb_counter_enable) = '1' then 
        analyzer_input_left_avalon_slave_arb_share_counter <= analyzer_input_left_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --analyzer_input_left_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      analyzer_input_left_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((analyzer_input_left_avalon_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_analyzer_input_left_avalon_slave)) OR ((end_xfer_arb_share_counter_term_analyzer_input_left_avalon_slave AND NOT analyzer_input_left_avalon_slave_non_bursting_master_requests)))) = '1' then 
        analyzer_input_left_avalon_slave_slavearbiterlockenable <= or_reduce(analyzer_input_left_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master analyzer_input_left/avalon_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= analyzer_input_left_avalon_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --analyzer_input_left_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  analyzer_input_left_avalon_slave_slavearbiterlockenable2 <= or_reduce(analyzer_input_left_avalon_slave_arb_share_counter_next_value);
  --cpu/data_master analyzer_input_left/avalon_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= analyzer_input_left_avalon_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --analyzer_input_left_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  analyzer_input_left_avalon_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_analyzer_input_left_avalon_slave <= internal_cpu_data_master_requests_analyzer_input_left_avalon_slave;
  --master is always granted when requested
  internal_cpu_data_master_granted_analyzer_input_left_avalon_slave <= internal_cpu_data_master_qualified_request_analyzer_input_left_avalon_slave;
  --cpu/data_master saved-grant analyzer_input_left/avalon_slave, which is an e_assign
  cpu_data_master_saved_grant_analyzer_input_left_avalon_slave <= internal_cpu_data_master_requests_analyzer_input_left_avalon_slave;
  --allow new arb cycle for analyzer_input_left/avalon_slave, which is an e_assign
  analyzer_input_left_avalon_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  analyzer_input_left_avalon_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  analyzer_input_left_avalon_slave_master_qreq_vector <= std_logic'('1');
  --analyzer_input_left_avalon_slave_reset_n assignment, which is an e_assign
  analyzer_input_left_avalon_slave_reset_n <= reset_n;
  --analyzer_input_left_avalon_slave_firsttransfer first transaction, which is an e_assign
  analyzer_input_left_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(analyzer_input_left_avalon_slave_begins_xfer) = '1'), analyzer_input_left_avalon_slave_unreg_firsttransfer, analyzer_input_left_avalon_slave_reg_firsttransfer);
  --analyzer_input_left_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  analyzer_input_left_avalon_slave_unreg_firsttransfer <= NOT ((analyzer_input_left_avalon_slave_slavearbiterlockenable AND analyzer_input_left_avalon_slave_any_continuerequest));
  --analyzer_input_left_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      analyzer_input_left_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(analyzer_input_left_avalon_slave_begins_xfer) = '1' then 
        analyzer_input_left_avalon_slave_reg_firsttransfer <= analyzer_input_left_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --analyzer_input_left_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  analyzer_input_left_avalon_slave_beginbursttransfer_internal <= analyzer_input_left_avalon_slave_begins_xfer;
  --analyzer_input_left_avalon_slave_read assignment, which is an e_mux
  analyzer_input_left_avalon_slave_read <= internal_cpu_data_master_granted_analyzer_input_left_avalon_slave AND cpu_data_master_read;
  shifted_address_to_analyzer_input_left_avalon_slave_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --d1_analyzer_input_left_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_analyzer_input_left_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_analyzer_input_left_avalon_slave_end_xfer <= analyzer_input_left_avalon_slave_end_xfer;
    end if;

  end process;

  --analyzer_input_left_avalon_slave_waits_for_read in a cycle, which is an e_mux
  analyzer_input_left_avalon_slave_waits_for_read <= analyzer_input_left_avalon_slave_in_a_read_cycle AND analyzer_input_left_avalon_slave_begins_xfer;
  --analyzer_input_left_avalon_slave_in_a_read_cycle assignment, which is an e_assign
  analyzer_input_left_avalon_slave_in_a_read_cycle <= internal_cpu_data_master_granted_analyzer_input_left_avalon_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= analyzer_input_left_avalon_slave_in_a_read_cycle;
  --analyzer_input_left_avalon_slave_waits_for_write in a cycle, which is an e_mux
  analyzer_input_left_avalon_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(analyzer_input_left_avalon_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --analyzer_input_left_avalon_slave_in_a_write_cycle assignment, which is an e_assign
  analyzer_input_left_avalon_slave_in_a_write_cycle <= internal_cpu_data_master_granted_analyzer_input_left_avalon_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= analyzer_input_left_avalon_slave_in_a_write_cycle;
  wait_for_analyzer_input_left_avalon_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_analyzer_input_left_avalon_slave <= internal_cpu_data_master_granted_analyzer_input_left_avalon_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_analyzer_input_left_avalon_slave <= internal_cpu_data_master_qualified_request_analyzer_input_left_avalon_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_analyzer_input_left_avalon_slave <= internal_cpu_data_master_requests_analyzer_input_left_avalon_slave;
--synthesis translate_off
    --analyzer_input_left/avalon_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity analyzer_input_right_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal analyzer_input_right_avalon_slave_readdata : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal analyzer_input_right_avalon_slave_read : OUT STD_LOGIC;
                 signal analyzer_input_right_avalon_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
                 signal analyzer_input_right_avalon_slave_reset_n : OUT STD_LOGIC;
                 signal cpu_data_master_granted_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                 signal d1_analyzer_input_right_avalon_slave_end_xfer : OUT STD_LOGIC
              );
end entity analyzer_input_right_avalon_slave_arbitrator;


architecture europa of analyzer_input_right_avalon_slave_arbitrator is
                signal analyzer_input_right_avalon_slave_allgrants :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal analyzer_input_right_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal analyzer_input_right_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal analyzer_input_right_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_begins_xfer :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_end_xfer :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_firsttransfer :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_grant_vector :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_in_a_read_cycle :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_in_a_write_cycle :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_master_qreq_vector :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_waits_for_read :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_waits_for_write :  STD_LOGIC;
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal shifted_address_to_analyzer_input_right_avalon_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_analyzer_input_right_avalon_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT analyzer_input_right_avalon_slave_end_xfer;
    end if;

  end process;

  analyzer_input_right_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_analyzer_input_right_avalon_slave);
  --assign analyzer_input_right_avalon_slave_readdata_from_sa = analyzer_input_right_avalon_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  analyzer_input_right_avalon_slave_readdata_from_sa <= analyzer_input_right_avalon_slave_readdata;
  internal_cpu_data_master_requests_analyzer_input_right_avalon_slave <= ((to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000110110000")))) AND ((cpu_data_master_read OR cpu_data_master_write)))) AND cpu_data_master_read;
  --analyzer_input_right_avalon_slave_arb_share_counter set values, which is an e_mux
  analyzer_input_right_avalon_slave_arb_share_set_values <= std_logic_vector'("001");
  --analyzer_input_right_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  analyzer_input_right_avalon_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_analyzer_input_right_avalon_slave;
  --analyzer_input_right_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  analyzer_input_right_avalon_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --analyzer_input_right_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  analyzer_input_right_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(analyzer_input_right_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (analyzer_input_right_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(analyzer_input_right_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (analyzer_input_right_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --analyzer_input_right_avalon_slave_allgrants all slave grants, which is an e_mux
  analyzer_input_right_avalon_slave_allgrants <= analyzer_input_right_avalon_slave_grant_vector;
  --analyzer_input_right_avalon_slave_end_xfer assignment, which is an e_assign
  analyzer_input_right_avalon_slave_end_xfer <= NOT ((analyzer_input_right_avalon_slave_waits_for_read OR analyzer_input_right_avalon_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_analyzer_input_right_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_analyzer_input_right_avalon_slave <= analyzer_input_right_avalon_slave_end_xfer AND (((NOT analyzer_input_right_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --analyzer_input_right_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  analyzer_input_right_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_analyzer_input_right_avalon_slave AND analyzer_input_right_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_analyzer_input_right_avalon_slave AND NOT analyzer_input_right_avalon_slave_non_bursting_master_requests));
  --analyzer_input_right_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      analyzer_input_right_avalon_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(analyzer_input_right_avalon_slave_arb_counter_enable) = '1' then 
        analyzer_input_right_avalon_slave_arb_share_counter <= analyzer_input_right_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --analyzer_input_right_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      analyzer_input_right_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((analyzer_input_right_avalon_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_analyzer_input_right_avalon_slave)) OR ((end_xfer_arb_share_counter_term_analyzer_input_right_avalon_slave AND NOT analyzer_input_right_avalon_slave_non_bursting_master_requests)))) = '1' then 
        analyzer_input_right_avalon_slave_slavearbiterlockenable <= or_reduce(analyzer_input_right_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master analyzer_input_right/avalon_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= analyzer_input_right_avalon_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --analyzer_input_right_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  analyzer_input_right_avalon_slave_slavearbiterlockenable2 <= or_reduce(analyzer_input_right_avalon_slave_arb_share_counter_next_value);
  --cpu/data_master analyzer_input_right/avalon_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= analyzer_input_right_avalon_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --analyzer_input_right_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  analyzer_input_right_avalon_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_analyzer_input_right_avalon_slave <= internal_cpu_data_master_requests_analyzer_input_right_avalon_slave;
  --master is always granted when requested
  internal_cpu_data_master_granted_analyzer_input_right_avalon_slave <= internal_cpu_data_master_qualified_request_analyzer_input_right_avalon_slave;
  --cpu/data_master saved-grant analyzer_input_right/avalon_slave, which is an e_assign
  cpu_data_master_saved_grant_analyzer_input_right_avalon_slave <= internal_cpu_data_master_requests_analyzer_input_right_avalon_slave;
  --allow new arb cycle for analyzer_input_right/avalon_slave, which is an e_assign
  analyzer_input_right_avalon_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  analyzer_input_right_avalon_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  analyzer_input_right_avalon_slave_master_qreq_vector <= std_logic'('1');
  --analyzer_input_right_avalon_slave_reset_n assignment, which is an e_assign
  analyzer_input_right_avalon_slave_reset_n <= reset_n;
  --analyzer_input_right_avalon_slave_firsttransfer first transaction, which is an e_assign
  analyzer_input_right_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(analyzer_input_right_avalon_slave_begins_xfer) = '1'), analyzer_input_right_avalon_slave_unreg_firsttransfer, analyzer_input_right_avalon_slave_reg_firsttransfer);
  --analyzer_input_right_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  analyzer_input_right_avalon_slave_unreg_firsttransfer <= NOT ((analyzer_input_right_avalon_slave_slavearbiterlockenable AND analyzer_input_right_avalon_slave_any_continuerequest));
  --analyzer_input_right_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      analyzer_input_right_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(analyzer_input_right_avalon_slave_begins_xfer) = '1' then 
        analyzer_input_right_avalon_slave_reg_firsttransfer <= analyzer_input_right_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --analyzer_input_right_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  analyzer_input_right_avalon_slave_beginbursttransfer_internal <= analyzer_input_right_avalon_slave_begins_xfer;
  --analyzer_input_right_avalon_slave_read assignment, which is an e_mux
  analyzer_input_right_avalon_slave_read <= internal_cpu_data_master_granted_analyzer_input_right_avalon_slave AND cpu_data_master_read;
  shifted_address_to_analyzer_input_right_avalon_slave_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --d1_analyzer_input_right_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_analyzer_input_right_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_analyzer_input_right_avalon_slave_end_xfer <= analyzer_input_right_avalon_slave_end_xfer;
    end if;

  end process;

  --analyzer_input_right_avalon_slave_waits_for_read in a cycle, which is an e_mux
  analyzer_input_right_avalon_slave_waits_for_read <= analyzer_input_right_avalon_slave_in_a_read_cycle AND analyzer_input_right_avalon_slave_begins_xfer;
  --analyzer_input_right_avalon_slave_in_a_read_cycle assignment, which is an e_assign
  analyzer_input_right_avalon_slave_in_a_read_cycle <= internal_cpu_data_master_granted_analyzer_input_right_avalon_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= analyzer_input_right_avalon_slave_in_a_read_cycle;
  --analyzer_input_right_avalon_slave_waits_for_write in a cycle, which is an e_mux
  analyzer_input_right_avalon_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(analyzer_input_right_avalon_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --analyzer_input_right_avalon_slave_in_a_write_cycle assignment, which is an e_assign
  analyzer_input_right_avalon_slave_in_a_write_cycle <= internal_cpu_data_master_granted_analyzer_input_right_avalon_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= analyzer_input_right_avalon_slave_in_a_write_cycle;
  wait_for_analyzer_input_right_avalon_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_analyzer_input_right_avalon_slave <= internal_cpu_data_master_granted_analyzer_input_right_avalon_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_analyzer_input_right_avalon_slave <= internal_cpu_data_master_qualified_request_analyzer_input_right_avalon_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_analyzer_input_right_avalon_slave <= internal_cpu_data_master_requests_analyzer_input_right_avalon_slave;
--synthesis translate_off
    --analyzer_input_right/avalon_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity audio_and_video_config_0_avalon_on_board_config_slave_arbitrator is 
        port (
              -- inputs:
                 signal audio_and_video_config_0_avalon_on_board_config_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal audio_and_video_config_0_avalon_on_board_config_slave_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal audio_and_video_config_0_avalon_on_board_config_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal audio_and_video_config_0_avalon_on_board_config_slave_chipselect : OUT STD_LOGIC;
                 signal audio_and_video_config_0_avalon_on_board_config_slave_read : OUT STD_LOGIC;
                 signal audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal audio_and_video_config_0_avalon_on_board_config_slave_reset : OUT STD_LOGIC;
                 signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal audio_and_video_config_0_avalon_on_board_config_slave_write : OUT STD_LOGIC;
                 signal audio_and_video_config_0_avalon_on_board_config_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                 signal d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC
              );
end entity audio_and_video_config_0_avalon_on_board_config_slave_arbitrator;


architecture europa of audio_and_video_config_0_avalon_on_board_config_slave_arbitrator is
                signal audio_and_video_config_0_avalon_on_board_config_slave_allgrants :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_any_continuerequest :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_arb_counter_enable :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal audio_and_video_config_0_avalon_on_board_config_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal audio_and_video_config_0_avalon_on_board_config_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_begins_xfer :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_end_xfer :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_firsttransfer :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_grant_vector :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_in_a_read_cycle :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_in_a_write_cycle :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_master_qreq_vector :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_non_bursting_master_requests :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_reg_firsttransfer :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_unreg_firsttransfer :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_waits_for_read :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_waits_for_write :  STD_LOGIC;
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_audio_and_video_config_0_avalon_on_board_config_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_audio_and_video_config_0_avalon_on_board_config_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT audio_and_video_config_0_avalon_on_board_config_slave_end_xfer;
    end if;

  end process;

  audio_and_video_config_0_avalon_on_board_config_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave);
  --assign audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa = audio_and_video_config_0_avalon_on_board_config_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa <= audio_and_video_config_0_avalon_on_board_config_slave_readdata;
  internal_cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("110100000011000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa = audio_and_video_config_0_avalon_on_board_config_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa <= audio_and_video_config_0_avalon_on_board_config_slave_waitrequest;
  --registered rdv signal_name registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave assignment, which is an e_assign
  registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave <= cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register_in;
  --audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter set values, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_arb_share_set_values <= std_logic_vector'("001");
  --audio_and_video_config_0_avalon_on_board_config_slave_non_bursting_master_requests mux, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave;
  --audio_and_video_config_0_avalon_on_board_config_slave_any_bursting_master_saved_grant mux, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter_next_value assignment, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(audio_and_video_config_0_avalon_on_board_config_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (audio_and_video_config_0_avalon_on_board_config_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --audio_and_video_config_0_avalon_on_board_config_slave_allgrants all slave grants, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_allgrants <= audio_and_video_config_0_avalon_on_board_config_slave_grant_vector;
  --audio_and_video_config_0_avalon_on_board_config_slave_end_xfer assignment, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_end_xfer <= NOT ((audio_and_video_config_0_avalon_on_board_config_slave_waits_for_read OR audio_and_video_config_0_avalon_on_board_config_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_audio_and_video_config_0_avalon_on_board_config_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_audio_and_video_config_0_avalon_on_board_config_slave <= audio_and_video_config_0_avalon_on_board_config_slave_end_xfer AND (((NOT audio_and_video_config_0_avalon_on_board_config_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter arbitration counter enable, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_audio_and_video_config_0_avalon_on_board_config_slave AND audio_and_video_config_0_avalon_on_board_config_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_audio_and_video_config_0_avalon_on_board_config_slave AND NOT audio_and_video_config_0_avalon_on_board_config_slave_non_bursting_master_requests));
  --audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(audio_and_video_config_0_avalon_on_board_config_slave_arb_counter_enable) = '1' then 
        audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter <= audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((audio_and_video_config_0_avalon_on_board_config_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_audio_and_video_config_0_avalon_on_board_config_slave)) OR ((end_xfer_arb_share_counter_term_audio_and_video_config_0_avalon_on_board_config_slave AND NOT audio_and_video_config_0_avalon_on_board_config_slave_non_bursting_master_requests)))) = '1' then 
        audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable <= or_reduce(audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master audio_and_video_config_0/avalon_on_board_config_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable2 <= or_reduce(audio_and_video_config_0_avalon_on_board_config_slave_arb_share_counter_next_value);
  --cpu/data_master audio_and_video_config_0/avalon_on_board_config_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --audio_and_video_config_0_avalon_on_board_config_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave <= internal_cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave AND NOT ((((cpu_data_master_read AND (cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register))) OR (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write))));
  --cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register_in <= ((internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave AND cpu_data_master_read) AND NOT audio_and_video_config_0_avalon_on_board_config_slave_waits_for_read) AND NOT (cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register);
  --shift register p1 cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register) & A_ToStdLogicVector(cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register_in)));
  --cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register <= p1_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave, which is an e_mux
  cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave <= cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave_shift_register;
  --audio_and_video_config_0_avalon_on_board_config_slave_writedata mux, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave <= internal_cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave;
  --cpu/data_master saved-grant audio_and_video_config_0/avalon_on_board_config_slave, which is an e_assign
  cpu_data_master_saved_grant_audio_and_video_config_0_avalon_on_board_config_slave <= internal_cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave;
  --allow new arb cycle for audio_and_video_config_0/avalon_on_board_config_slave, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  audio_and_video_config_0_avalon_on_board_config_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  audio_and_video_config_0_avalon_on_board_config_slave_master_qreq_vector <= std_logic'('1');
  --~audio_and_video_config_0_avalon_on_board_config_slave_reset assignment, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_reset <= NOT reset_n;
  audio_and_video_config_0_avalon_on_board_config_slave_chipselect <= internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave;
  --audio_and_video_config_0_avalon_on_board_config_slave_firsttransfer first transaction, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_firsttransfer <= A_WE_StdLogic((std_logic'(audio_and_video_config_0_avalon_on_board_config_slave_begins_xfer) = '1'), audio_and_video_config_0_avalon_on_board_config_slave_unreg_firsttransfer, audio_and_video_config_0_avalon_on_board_config_slave_reg_firsttransfer);
  --audio_and_video_config_0_avalon_on_board_config_slave_unreg_firsttransfer first transaction, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_unreg_firsttransfer <= NOT ((audio_and_video_config_0_avalon_on_board_config_slave_slavearbiterlockenable AND audio_and_video_config_0_avalon_on_board_config_slave_any_continuerequest));
  --audio_and_video_config_0_avalon_on_board_config_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      audio_and_video_config_0_avalon_on_board_config_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(audio_and_video_config_0_avalon_on_board_config_slave_begins_xfer) = '1' then 
        audio_and_video_config_0_avalon_on_board_config_slave_reg_firsttransfer <= audio_and_video_config_0_avalon_on_board_config_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --audio_and_video_config_0_avalon_on_board_config_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_beginbursttransfer_internal <= audio_and_video_config_0_avalon_on_board_config_slave_begins_xfer;
  --audio_and_video_config_0_avalon_on_board_config_slave_read assignment, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_read <= internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave AND cpu_data_master_read;
  --audio_and_video_config_0_avalon_on_board_config_slave_write assignment, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_write <= internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave AND cpu_data_master_write;
  shifted_address_to_audio_and_video_config_0_avalon_on_board_config_slave_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --audio_and_video_config_0_avalon_on_board_config_slave_address mux, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_address <= A_EXT (A_SRL(shifted_address_to_audio_and_video_config_0_avalon_on_board_config_slave_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer <= audio_and_video_config_0_avalon_on_board_config_slave_end_xfer;
    end if;

  end process;

  --audio_and_video_config_0_avalon_on_board_config_slave_waits_for_read in a cycle, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_waits_for_read <= audio_and_video_config_0_avalon_on_board_config_slave_in_a_read_cycle AND internal_audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa;
  --audio_and_video_config_0_avalon_on_board_config_slave_in_a_read_cycle assignment, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_in_a_read_cycle <= internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= audio_and_video_config_0_avalon_on_board_config_slave_in_a_read_cycle;
  --audio_and_video_config_0_avalon_on_board_config_slave_waits_for_write in a cycle, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_waits_for_write <= audio_and_video_config_0_avalon_on_board_config_slave_in_a_write_cycle AND internal_audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa;
  --audio_and_video_config_0_avalon_on_board_config_slave_in_a_write_cycle assignment, which is an e_assign
  audio_and_video_config_0_avalon_on_board_config_slave_in_a_write_cycle <= internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= audio_and_video_config_0_avalon_on_board_config_slave_in_a_write_cycle;
  wait_for_audio_and_video_config_0_avalon_on_board_config_slave_counter <= std_logic'('0');
  --audio_and_video_config_0_avalon_on_board_config_slave_byteenable byte enable port mux, which is an e_mux
  audio_and_video_config_0_avalon_on_board_config_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa <= internal_audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave <= internal_cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave <= internal_cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave <= internal_cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave;
--synthesis translate_off
    --audio_and_video_config_0/avalon_on_board_config_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity character_buffer_avalon_char_buffer_slave_arbitrator is 
        port (
              -- inputs:
                 signal character_buffer_avalon_char_buffer_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal character_buffer_avalon_char_buffer_slave_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal character_buffer_avalon_char_buffer_slave_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal character_buffer_avalon_char_buffer_slave_chipselect : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_buffer_slave_read : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_buffer_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal character_buffer_avalon_char_buffer_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_buffer_slave_write : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_buffer_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal cpu_data_master_granted_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                 signal d1_character_buffer_avalon_char_buffer_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC
              );
end entity character_buffer_avalon_char_buffer_slave_arbitrator;


architecture europa of character_buffer_avalon_char_buffer_slave_arbitrator is
                signal character_buffer_avalon_char_buffer_slave_allgrants :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_any_continuerequest :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_arb_counter_enable :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal character_buffer_avalon_char_buffer_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal character_buffer_avalon_char_buffer_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal character_buffer_avalon_char_buffer_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_begins_xfer :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_end_xfer :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_firsttransfer :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_grant_vector :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_in_a_read_cycle :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_in_a_write_cycle :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_master_qreq_vector :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_non_bursting_master_requests :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_pretend_byte_enable :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_reg_firsttransfer :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_slavearbiterlockenable :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_unreg_firsttransfer :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_waits_for_read :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_waits_for_write :  STD_LOGIC;
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_0 :  STD_LOGIC;
                signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_1 :  STD_LOGIC;
                signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_3 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_character_buffer_avalon_char_buffer_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register :  STD_LOGIC;
                signal wait_for_character_buffer_avalon_char_buffer_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT character_buffer_avalon_char_buffer_slave_end_xfer;
    end if;

  end process;

  character_buffer_avalon_char_buffer_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave);
  --assign character_buffer_avalon_char_buffer_slave_readdata_from_sa = character_buffer_avalon_char_buffer_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  character_buffer_avalon_char_buffer_slave_readdata_from_sa <= character_buffer_avalon_char_buffer_slave_readdata;
  internal_cpu_data_master_requests_character_buffer_avalon_char_buffer_slave <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("110100000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign character_buffer_avalon_char_buffer_slave_waitrequest_from_sa = character_buffer_avalon_char_buffer_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_character_buffer_avalon_char_buffer_slave_waitrequest_from_sa <= character_buffer_avalon_char_buffer_slave_waitrequest;
  --registered rdv signal_name registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave assignment, which is an e_assign
  registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave <= cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register_in;
  --character_buffer_avalon_char_buffer_slave_arb_share_counter set values, which is an e_mux
  character_buffer_avalon_char_buffer_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000001")), 3);
  --character_buffer_avalon_char_buffer_slave_non_bursting_master_requests mux, which is an e_mux
  character_buffer_avalon_char_buffer_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_character_buffer_avalon_char_buffer_slave;
  --character_buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant mux, which is an e_mux
  character_buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --character_buffer_avalon_char_buffer_slave_arb_share_counter_next_value assignment, which is an e_assign
  character_buffer_avalon_char_buffer_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(character_buffer_avalon_char_buffer_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (character_buffer_avalon_char_buffer_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(character_buffer_avalon_char_buffer_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (character_buffer_avalon_char_buffer_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --character_buffer_avalon_char_buffer_slave_allgrants all slave grants, which is an e_mux
  character_buffer_avalon_char_buffer_slave_allgrants <= character_buffer_avalon_char_buffer_slave_grant_vector;
  --character_buffer_avalon_char_buffer_slave_end_xfer assignment, which is an e_assign
  character_buffer_avalon_char_buffer_slave_end_xfer <= NOT ((character_buffer_avalon_char_buffer_slave_waits_for_read OR character_buffer_avalon_char_buffer_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_character_buffer_avalon_char_buffer_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_character_buffer_avalon_char_buffer_slave <= character_buffer_avalon_char_buffer_slave_end_xfer AND (((NOT character_buffer_avalon_char_buffer_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --character_buffer_avalon_char_buffer_slave_arb_share_counter arbitration counter enable, which is an e_assign
  character_buffer_avalon_char_buffer_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_character_buffer_avalon_char_buffer_slave AND character_buffer_avalon_char_buffer_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_character_buffer_avalon_char_buffer_slave AND NOT character_buffer_avalon_char_buffer_slave_non_bursting_master_requests));
  --character_buffer_avalon_char_buffer_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      character_buffer_avalon_char_buffer_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(character_buffer_avalon_char_buffer_slave_arb_counter_enable) = '1' then 
        character_buffer_avalon_char_buffer_slave_arb_share_counter <= character_buffer_avalon_char_buffer_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --character_buffer_avalon_char_buffer_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      character_buffer_avalon_char_buffer_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((character_buffer_avalon_char_buffer_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_character_buffer_avalon_char_buffer_slave)) OR ((end_xfer_arb_share_counter_term_character_buffer_avalon_char_buffer_slave AND NOT character_buffer_avalon_char_buffer_slave_non_bursting_master_requests)))) = '1' then 
        character_buffer_avalon_char_buffer_slave_slavearbiterlockenable <= or_reduce(character_buffer_avalon_char_buffer_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master character_buffer/avalon_char_buffer_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= character_buffer_avalon_char_buffer_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --character_buffer_avalon_char_buffer_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  character_buffer_avalon_char_buffer_slave_slavearbiterlockenable2 <= or_reduce(character_buffer_avalon_char_buffer_slave_arb_share_counter_next_value);
  --cpu/data_master character_buffer/avalon_char_buffer_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= character_buffer_avalon_char_buffer_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --character_buffer_avalon_char_buffer_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  character_buffer_avalon_char_buffer_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave <= internal_cpu_data_master_requests_character_buffer_avalon_char_buffer_slave AND NOT ((((cpu_data_master_read AND (cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register))) OR (((((NOT cpu_data_master_waitrequest OR cpu_data_master_no_byte_enables_and_last_term) OR NOT(internal_cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave))) AND cpu_data_master_write))));
  --cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register_in <= ((internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave AND cpu_data_master_read) AND NOT character_buffer_avalon_char_buffer_slave_waits_for_read) AND NOT (cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register);
  --shift register p1 cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register) & A_ToStdLogicVector(cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register_in)));
  --cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register <= p1_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave, which is an e_mux
  cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave <= cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave_shift_register;
  --character_buffer_avalon_char_buffer_slave_writedata mux, which is an e_mux
  character_buffer_avalon_char_buffer_slave_writedata <= cpu_data_master_dbs_write_8;
  --master is always granted when requested
  internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave <= internal_cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave;
  --cpu/data_master saved-grant character_buffer/avalon_char_buffer_slave, which is an e_assign
  cpu_data_master_saved_grant_character_buffer_avalon_char_buffer_slave <= internal_cpu_data_master_requests_character_buffer_avalon_char_buffer_slave;
  --allow new arb cycle for character_buffer/avalon_char_buffer_slave, which is an e_assign
  character_buffer_avalon_char_buffer_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  character_buffer_avalon_char_buffer_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  character_buffer_avalon_char_buffer_slave_master_qreq_vector <= std_logic'('1');
  character_buffer_avalon_char_buffer_slave_chipselect <= internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave;
  --character_buffer_avalon_char_buffer_slave_firsttransfer first transaction, which is an e_assign
  character_buffer_avalon_char_buffer_slave_firsttransfer <= A_WE_StdLogic((std_logic'(character_buffer_avalon_char_buffer_slave_begins_xfer) = '1'), character_buffer_avalon_char_buffer_slave_unreg_firsttransfer, character_buffer_avalon_char_buffer_slave_reg_firsttransfer);
  --character_buffer_avalon_char_buffer_slave_unreg_firsttransfer first transaction, which is an e_assign
  character_buffer_avalon_char_buffer_slave_unreg_firsttransfer <= NOT ((character_buffer_avalon_char_buffer_slave_slavearbiterlockenable AND character_buffer_avalon_char_buffer_slave_any_continuerequest));
  --character_buffer_avalon_char_buffer_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      character_buffer_avalon_char_buffer_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(character_buffer_avalon_char_buffer_slave_begins_xfer) = '1' then 
        character_buffer_avalon_char_buffer_slave_reg_firsttransfer <= character_buffer_avalon_char_buffer_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --character_buffer_avalon_char_buffer_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  character_buffer_avalon_char_buffer_slave_beginbursttransfer_internal <= character_buffer_avalon_char_buffer_slave_begins_xfer;
  --character_buffer_avalon_char_buffer_slave_read assignment, which is an e_mux
  character_buffer_avalon_char_buffer_slave_read <= internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave AND cpu_data_master_read;
  --character_buffer_avalon_char_buffer_slave_write assignment, which is an e_mux
  character_buffer_avalon_char_buffer_slave_write <= ((internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave AND cpu_data_master_write)) AND character_buffer_avalon_char_buffer_slave_pretend_byte_enable;
  --character_buffer_avalon_char_buffer_slave_address mux, which is an e_mux
  character_buffer_avalon_char_buffer_slave_address <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & cpu_data_master_dbs_address(1 DOWNTO 0)), 13);
  --d1_character_buffer_avalon_char_buffer_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_character_buffer_avalon_char_buffer_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_character_buffer_avalon_char_buffer_slave_end_xfer <= character_buffer_avalon_char_buffer_slave_end_xfer;
    end if;

  end process;

  --character_buffer_avalon_char_buffer_slave_waits_for_read in a cycle, which is an e_mux
  character_buffer_avalon_char_buffer_slave_waits_for_read <= character_buffer_avalon_char_buffer_slave_in_a_read_cycle AND internal_character_buffer_avalon_char_buffer_slave_waitrequest_from_sa;
  --character_buffer_avalon_char_buffer_slave_in_a_read_cycle assignment, which is an e_assign
  character_buffer_avalon_char_buffer_slave_in_a_read_cycle <= internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= character_buffer_avalon_char_buffer_slave_in_a_read_cycle;
  --character_buffer_avalon_char_buffer_slave_waits_for_write in a cycle, which is an e_mux
  character_buffer_avalon_char_buffer_slave_waits_for_write <= character_buffer_avalon_char_buffer_slave_in_a_write_cycle AND internal_character_buffer_avalon_char_buffer_slave_waitrequest_from_sa;
  --character_buffer_avalon_char_buffer_slave_in_a_write_cycle assignment, which is an e_assign
  character_buffer_avalon_char_buffer_slave_in_a_write_cycle <= internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= character_buffer_avalon_char_buffer_slave_in_a_write_cycle;
  wait_for_character_buffer_avalon_char_buffer_slave_counter <= std_logic'('0');
  --character_buffer_avalon_char_buffer_slave_pretend_byte_enable byte enable port mux, which is an e_mux
  character_buffer_avalon_char_buffer_slave_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  (cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_3, cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_2, cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_1, cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_0) <= cpu_data_master_byteenable;
  internal_cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave <= A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_0, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_1, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_2, cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave_segment_3)));
  --vhdl renameroo for output signals
  character_buffer_avalon_char_buffer_slave_waitrequest_from_sa <= internal_character_buffer_avalon_char_buffer_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave <= internal_cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave;
  --vhdl renameroo for output signals
  cpu_data_master_granted_character_buffer_avalon_char_buffer_slave <= internal_cpu_data_master_granted_character_buffer_avalon_char_buffer_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave <= internal_cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_character_buffer_avalon_char_buffer_slave <= internal_cpu_data_master_requests_character_buffer_avalon_char_buffer_slave;
--synthesis translate_off
    --character_buffer/avalon_char_buffer_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity character_buffer_avalon_char_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal character_buffer_avalon_char_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal character_buffer_avalon_char_control_slave_address : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_control_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal character_buffer_avalon_char_control_slave_chipselect : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_control_slave_read : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal character_buffer_avalon_char_control_slave_reset : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_control_slave_write : OUT STD_LOGIC;
                 signal character_buffer_avalon_char_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_granted_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                 signal d1_character_buffer_avalon_char_control_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : OUT STD_LOGIC
              );
end entity character_buffer_avalon_char_control_slave_arbitrator;


architecture europa of character_buffer_avalon_char_control_slave_arbitrator is
                signal character_buffer_avalon_char_control_slave_allgrants :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_any_continuerequest :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_arb_counter_enable :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal character_buffer_avalon_char_control_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal character_buffer_avalon_char_control_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal character_buffer_avalon_char_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_begins_xfer :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_end_xfer :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_firsttransfer :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_grant_vector :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_master_qreq_vector :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_waits_for_read :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_waits_for_write :  STD_LOGIC;
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register :  STD_LOGIC;
                signal shifted_address_to_character_buffer_avalon_char_control_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_character_buffer_avalon_char_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT character_buffer_avalon_char_control_slave_end_xfer;
    end if;

  end process;

  character_buffer_avalon_char_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave);
  --assign character_buffer_avalon_char_control_slave_readdata_from_sa = character_buffer_avalon_char_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  character_buffer_avalon_char_control_slave_readdata_from_sa <= character_buffer_avalon_char_control_slave_readdata;
  internal_cpu_data_master_requests_character_buffer_avalon_char_control_slave <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("110100000011000111100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --registered rdv signal_name registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave assignment, which is an e_assign
  registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave <= cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register_in;
  --character_buffer_avalon_char_control_slave_arb_share_counter set values, which is an e_mux
  character_buffer_avalon_char_control_slave_arb_share_set_values <= std_logic_vector'("001");
  --character_buffer_avalon_char_control_slave_non_bursting_master_requests mux, which is an e_mux
  character_buffer_avalon_char_control_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_character_buffer_avalon_char_control_slave;
  --character_buffer_avalon_char_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  character_buffer_avalon_char_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --character_buffer_avalon_char_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  character_buffer_avalon_char_control_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(character_buffer_avalon_char_control_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (character_buffer_avalon_char_control_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(character_buffer_avalon_char_control_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (character_buffer_avalon_char_control_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --character_buffer_avalon_char_control_slave_allgrants all slave grants, which is an e_mux
  character_buffer_avalon_char_control_slave_allgrants <= character_buffer_avalon_char_control_slave_grant_vector;
  --character_buffer_avalon_char_control_slave_end_xfer assignment, which is an e_assign
  character_buffer_avalon_char_control_slave_end_xfer <= NOT ((character_buffer_avalon_char_control_slave_waits_for_read OR character_buffer_avalon_char_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_character_buffer_avalon_char_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_character_buffer_avalon_char_control_slave <= character_buffer_avalon_char_control_slave_end_xfer AND (((NOT character_buffer_avalon_char_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --character_buffer_avalon_char_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  character_buffer_avalon_char_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_character_buffer_avalon_char_control_slave AND character_buffer_avalon_char_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_character_buffer_avalon_char_control_slave AND NOT character_buffer_avalon_char_control_slave_non_bursting_master_requests));
  --character_buffer_avalon_char_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      character_buffer_avalon_char_control_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(character_buffer_avalon_char_control_slave_arb_counter_enable) = '1' then 
        character_buffer_avalon_char_control_slave_arb_share_counter <= character_buffer_avalon_char_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --character_buffer_avalon_char_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      character_buffer_avalon_char_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((character_buffer_avalon_char_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_character_buffer_avalon_char_control_slave)) OR ((end_xfer_arb_share_counter_term_character_buffer_avalon_char_control_slave AND NOT character_buffer_avalon_char_control_slave_non_bursting_master_requests)))) = '1' then 
        character_buffer_avalon_char_control_slave_slavearbiterlockenable <= or_reduce(character_buffer_avalon_char_control_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master character_buffer/avalon_char_control_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= character_buffer_avalon_char_control_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --character_buffer_avalon_char_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  character_buffer_avalon_char_control_slave_slavearbiterlockenable2 <= or_reduce(character_buffer_avalon_char_control_slave_arb_share_counter_next_value);
  --cpu/data_master character_buffer/avalon_char_control_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= character_buffer_avalon_char_control_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --character_buffer_avalon_char_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  character_buffer_avalon_char_control_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave <= internal_cpu_data_master_requests_character_buffer_avalon_char_control_slave AND NOT ((((cpu_data_master_read AND (cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register))) OR (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write))));
  --cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register_in <= ((internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave AND cpu_data_master_read) AND NOT character_buffer_avalon_char_control_slave_waits_for_read) AND NOT (cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register);
  --shift register p1 cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register) & A_ToStdLogicVector(cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register_in)));
  --cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register <= p1_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave, which is an e_mux
  cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave <= cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave_shift_register;
  --character_buffer_avalon_char_control_slave_writedata mux, which is an e_mux
  character_buffer_avalon_char_control_slave_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave <= internal_cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave;
  --cpu/data_master saved-grant character_buffer/avalon_char_control_slave, which is an e_assign
  cpu_data_master_saved_grant_character_buffer_avalon_char_control_slave <= internal_cpu_data_master_requests_character_buffer_avalon_char_control_slave;
  --allow new arb cycle for character_buffer/avalon_char_control_slave, which is an e_assign
  character_buffer_avalon_char_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  character_buffer_avalon_char_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  character_buffer_avalon_char_control_slave_master_qreq_vector <= std_logic'('1');
  --~character_buffer_avalon_char_control_slave_reset assignment, which is an e_assign
  character_buffer_avalon_char_control_slave_reset <= NOT reset_n;
  character_buffer_avalon_char_control_slave_chipselect <= internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave;
  --character_buffer_avalon_char_control_slave_firsttransfer first transaction, which is an e_assign
  character_buffer_avalon_char_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(character_buffer_avalon_char_control_slave_begins_xfer) = '1'), character_buffer_avalon_char_control_slave_unreg_firsttransfer, character_buffer_avalon_char_control_slave_reg_firsttransfer);
  --character_buffer_avalon_char_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  character_buffer_avalon_char_control_slave_unreg_firsttransfer <= NOT ((character_buffer_avalon_char_control_slave_slavearbiterlockenable AND character_buffer_avalon_char_control_slave_any_continuerequest));
  --character_buffer_avalon_char_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      character_buffer_avalon_char_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(character_buffer_avalon_char_control_slave_begins_xfer) = '1' then 
        character_buffer_avalon_char_control_slave_reg_firsttransfer <= character_buffer_avalon_char_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --character_buffer_avalon_char_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  character_buffer_avalon_char_control_slave_beginbursttransfer_internal <= character_buffer_avalon_char_control_slave_begins_xfer;
  --character_buffer_avalon_char_control_slave_read assignment, which is an e_mux
  character_buffer_avalon_char_control_slave_read <= internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave AND cpu_data_master_read;
  --character_buffer_avalon_char_control_slave_write assignment, which is an e_mux
  character_buffer_avalon_char_control_slave_write <= internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave AND cpu_data_master_write;
  shifted_address_to_character_buffer_avalon_char_control_slave_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --character_buffer_avalon_char_control_slave_address mux, which is an e_mux
  character_buffer_avalon_char_control_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_character_buffer_avalon_char_control_slave_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_character_buffer_avalon_char_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_character_buffer_avalon_char_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_character_buffer_avalon_char_control_slave_end_xfer <= character_buffer_avalon_char_control_slave_end_xfer;
    end if;

  end process;

  --character_buffer_avalon_char_control_slave_waits_for_read in a cycle, which is an e_mux
  character_buffer_avalon_char_control_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(character_buffer_avalon_char_control_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --character_buffer_avalon_char_control_slave_in_a_read_cycle assignment, which is an e_assign
  character_buffer_avalon_char_control_slave_in_a_read_cycle <= internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= character_buffer_avalon_char_control_slave_in_a_read_cycle;
  --character_buffer_avalon_char_control_slave_waits_for_write in a cycle, which is an e_mux
  character_buffer_avalon_char_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(character_buffer_avalon_char_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --character_buffer_avalon_char_control_slave_in_a_write_cycle assignment, which is an e_assign
  character_buffer_avalon_char_control_slave_in_a_write_cycle <= internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= character_buffer_avalon_char_control_slave_in_a_write_cycle;
  wait_for_character_buffer_avalon_char_control_slave_counter <= std_logic'('0');
  --character_buffer_avalon_char_control_slave_byteenable byte enable port mux, which is an e_mux
  character_buffer_avalon_char_control_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_data_master_granted_character_buffer_avalon_char_control_slave <= internal_cpu_data_master_granted_character_buffer_avalon_char_control_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave <= internal_cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_character_buffer_avalon_char_control_slave <= internal_cpu_data_master_requests_character_buffer_avalon_char_control_slave;
--synthesis translate_off
    --character_buffer/avalon_char_control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity character_buffer_avalon_char_source_arbitrator is 
        port (
              -- inputs:
                 signal alpha_blending_avalon_foreground_sink_ready_from_sa : IN STD_LOGIC;
                 signal character_buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                 signal character_buffer_avalon_char_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal character_buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                 signal character_buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                 signal character_buffer_avalon_char_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal character_buffer_avalon_char_source_ready : OUT STD_LOGIC
              );
end entity character_buffer_avalon_char_source_arbitrator;


architecture europa of character_buffer_avalon_char_source_arbitrator is

begin

  --mux character_buffer_avalon_char_source_ready, which is an e_mux
  character_buffer_avalon_char_source_ready <= alpha_blending_avalon_foreground_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_data_master_requests_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_instruction_master_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_write : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC
              );
end entity cpu_jtag_debug_module_arbitrator;


architecture europa of cpu_jtag_debug_module_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_jtag_debug_module_allgrants :  STD_LOGIC;
                signal cpu_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpu_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal cpu_jtag_debug_module_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal cpu_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal cpu_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal cpu_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal cpu_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpu_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal cpu_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpu_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_data_master_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_cpu_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  cpu_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_data_master_qualified_request_cpu_jtag_debug_module OR internal_cpu_instruction_master_qualified_request_cpu_jtag_debug_module));
  --assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_jtag_debug_module_readdata_from_sa <= cpu_jtag_debug_module_readdata;
  internal_cpu_data_master_requests_cpu_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("110100000010100000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  cpu_jtag_debug_module_arb_share_set_values <= std_logic_vector'("001");
  --cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  cpu_jtag_debug_module_non_bursting_master_requests <= ((internal_cpu_data_master_requests_cpu_jtag_debug_module OR internal_cpu_instruction_master_requests_cpu_jtag_debug_module) OR internal_cpu_data_master_requests_cpu_jtag_debug_module) OR internal_cpu_instruction_master_requests_cpu_jtag_debug_module;
  --cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  cpu_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  cpu_jtag_debug_module_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(cpu_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (cpu_jtag_debug_module_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(cpu_jtag_debug_module_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (cpu_jtag_debug_module_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  cpu_jtag_debug_module_allgrants <= (((or_reduce(cpu_jtag_debug_module_grant_vector)) OR (or_reduce(cpu_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_jtag_debug_module_grant_vector));
  --cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  cpu_jtag_debug_module_end_xfer <= NOT ((cpu_jtag_debug_module_waits_for_read OR cpu_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpu_jtag_debug_module <= cpu_jtag_debug_module_end_xfer AND (((NOT cpu_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  cpu_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND cpu_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND NOT cpu_jtag_debug_module_non_bursting_master_requests));
  --cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_arb_counter_enable) = '1' then 
        cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(cpu_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_cpu_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND NOT cpu_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        cpu_jtag_debug_module_slavearbiterlockenable <= or_reduce(cpu_jtag_debug_module_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= cpu_jtag_debug_module_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpu_jtag_debug_module_slavearbiterlockenable2 <= or_reduce(cpu_jtag_debug_module_arb_share_counter_next_value);
  --cpu/data_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= cpu_jtag_debug_module_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --cpu/instruction_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= cpu_jtag_debug_module_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= cpu_jtag_debug_module_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master granted cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_instruction_master_saved_grant_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpu_instruction_master_requests_cpu_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module))))));
    end if;

  end process;

  --cpu_instruction_master_continuerequest continued request, which is an e_mux
  cpu_instruction_master_continuerequest <= last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module AND internal_cpu_instruction_master_requests_cpu_jtag_debug_module;
  --cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  cpu_jtag_debug_module_any_continuerequest <= cpu_instruction_master_continuerequest OR cpu_data_master_continuerequest;
  internal_cpu_data_master_qualified_request_cpu_jtag_debug_module <= internal_cpu_data_master_requests_cpu_jtag_debug_module AND NOT (((((NOT cpu_data_master_waitrequest) AND cpu_data_master_write)) OR cpu_instruction_master_arbiterlock));
  --cpu_jtag_debug_module_writedata mux, which is an e_mux
  cpu_jtag_debug_module_writedata <= cpu_data_master_writedata;
  internal_cpu_instruction_master_requests_cpu_jtag_debug_module <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(23 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("110100000010100000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --cpu/data_master granted cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_data_master_saved_grant_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpu_data_master_requests_cpu_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module))))));
    end if;

  end process;

  --cpu_data_master_continuerequest continued request, which is an e_mux
  cpu_data_master_continuerequest <= last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module AND internal_cpu_data_master_requests_cpu_jtag_debug_module;
  internal_cpu_instruction_master_qualified_request_cpu_jtag_debug_module <= internal_cpu_instruction_master_requests_cpu_jtag_debug_module AND NOT ((((cpu_instruction_master_read AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (cpu_instruction_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000")))))) OR cpu_data_master_arbiterlock));
  --local readdatavalid cpu_instruction_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  cpu_instruction_master_read_data_valid_cpu_jtag_debug_module <= (internal_cpu_instruction_master_granted_cpu_jtag_debug_module AND cpu_instruction_master_read) AND NOT cpu_jtag_debug_module_waits_for_read;
  --allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  cpu_jtag_debug_module_allow_new_arb_cycle <= NOT cpu_data_master_arbiterlock AND NOT cpu_instruction_master_arbiterlock;
  --cpu/instruction_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  cpu_jtag_debug_module_master_qreq_vector(0) <= internal_cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  --cpu/instruction_master grant cpu/jtag_debug_module, which is an e_assign
  internal_cpu_instruction_master_granted_cpu_jtag_debug_module <= cpu_jtag_debug_module_grant_vector(0);
  --cpu/instruction_master saved-grant cpu/jtag_debug_module, which is an e_assign
  cpu_instruction_master_saved_grant_cpu_jtag_debug_module <= cpu_jtag_debug_module_arb_winner(0) AND internal_cpu_instruction_master_requests_cpu_jtag_debug_module;
  --cpu/data_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  cpu_jtag_debug_module_master_qreq_vector(1) <= internal_cpu_data_master_qualified_request_cpu_jtag_debug_module;
  --cpu/data_master grant cpu/jtag_debug_module, which is an e_assign
  internal_cpu_data_master_granted_cpu_jtag_debug_module <= cpu_jtag_debug_module_grant_vector(1);
  --cpu/data_master saved-grant cpu/jtag_debug_module, which is an e_assign
  cpu_data_master_saved_grant_cpu_jtag_debug_module <= cpu_jtag_debug_module_arb_winner(1) AND internal_cpu_data_master_requests_cpu_jtag_debug_module;
  --cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  cpu_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((cpu_jtag_debug_module_master_qreq_vector & cpu_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT cpu_jtag_debug_module_master_qreq_vector & NOT cpu_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (cpu_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  cpu_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((cpu_jtag_debug_module_allow_new_arb_cycle AND or_reduce(cpu_jtag_debug_module_grant_vector)))) = '1'), cpu_jtag_debug_module_grant_vector, cpu_jtag_debug_module_saved_chosen_master_vector);
  --saved cpu_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        cpu_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(cpu_jtag_debug_module_grant_vector)) = '1'), cpu_jtag_debug_module_grant_vector, cpu_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  cpu_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((cpu_jtag_debug_module_chosen_master_double_vector(1) OR cpu_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((cpu_jtag_debug_module_chosen_master_double_vector(0) OR cpu_jtag_debug_module_chosen_master_double_vector(2)))));
  --cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  cpu_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --cpu/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(cpu_jtag_debug_module_grant_vector)) = '1' then 
        cpu_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(cpu_jtag_debug_module_end_xfer) = '1'), cpu_jtag_debug_module_chosen_master_rot_left, cpu_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  cpu_jtag_debug_module_begintransfer <= cpu_jtag_debug_module_begins_xfer;
  --assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_jtag_debug_module_resetrequest_from_sa <= cpu_jtag_debug_module_resetrequest;
  cpu_jtag_debug_module_chipselect <= internal_cpu_data_master_granted_cpu_jtag_debug_module OR internal_cpu_instruction_master_granted_cpu_jtag_debug_module;
  --cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  cpu_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(cpu_jtag_debug_module_begins_xfer) = '1'), cpu_jtag_debug_module_unreg_firsttransfer, cpu_jtag_debug_module_reg_firsttransfer);
  --cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  cpu_jtag_debug_module_unreg_firsttransfer <= NOT ((cpu_jtag_debug_module_slavearbiterlockenable AND cpu_jtag_debug_module_any_continuerequest));
  --cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_begins_xfer) = '1' then 
        cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpu_jtag_debug_module_beginbursttransfer_internal <= cpu_jtag_debug_module_begins_xfer;
  --cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  cpu_jtag_debug_module_arbitration_holdoff_internal <= cpu_jtag_debug_module_begins_xfer AND cpu_jtag_debug_module_firsttransfer;
  --cpu_jtag_debug_module_write assignment, which is an e_mux
  cpu_jtag_debug_module_write <= internal_cpu_data_master_granted_cpu_jtag_debug_module AND cpu_data_master_write;
  shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --cpu_jtag_debug_module_address mux, which is an e_mux
  cpu_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_cpu_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master <= cpu_instruction_master_address_to_slave;
  --d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpu_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  --cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  cpu_jtag_debug_module_waits_for_read <= cpu_jtag_debug_module_in_a_read_cycle AND cpu_jtag_debug_module_begins_xfer;
  --cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  cpu_jtag_debug_module_in_a_read_cycle <= ((internal_cpu_data_master_granted_cpu_jtag_debug_module AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_cpu_jtag_debug_module AND cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpu_jtag_debug_module_in_a_read_cycle;
  --cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  cpu_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  cpu_jtag_debug_module_in_a_write_cycle <= internal_cpu_data_master_granted_cpu_jtag_debug_module AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpu_jtag_debug_module_in_a_write_cycle;
  wait_for_cpu_jtag_debug_module_counter <= std_logic'('0');
  --cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  cpu_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  cpu_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_cpu_jtag_debug_module <= internal_cpu_data_master_granted_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_cpu_jtag_debug_module <= internal_cpu_data_master_qualified_request_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_data_master_requests_cpu_jtag_debug_module <= internal_cpu_data_master_requests_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_cpu_jtag_debug_module <= internal_cpu_instruction_master_granted_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_cpu_jtag_debug_module <= internal_cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_cpu_jtag_debug_module <= internal_cpu_instruction_master_requests_cpu_jtag_debug_module;
--synthesis translate_off
    --cpu/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_granted_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_instruction_master_granted_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_data_master_saved_grant_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_saved_grant_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpu_custom_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_custom_instruction_master_multi_start : IN STD_LOGIC;
                 signal cpu_fpoint_s1_done_from_sa : IN STD_LOGIC;
                 signal cpu_fpoint_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_custom_instruction_master_multi_done : OUT STD_LOGIC;
                 signal cpu_custom_instruction_master_multi_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_custom_instruction_master_reset_n : OUT STD_LOGIC;
                 signal cpu_custom_instruction_master_start_cpu_fpoint_s1 : OUT STD_LOGIC;
                 signal cpu_fpoint_s1_select : OUT STD_LOGIC
              );
end entity cpu_custom_instruction_master_arbitrator;


architecture europa of cpu_custom_instruction_master_arbitrator is
                signal internal_cpu_fpoint_s1_select :  STD_LOGIC;

begin

  internal_cpu_fpoint_s1_select <= std_logic'('1');
  cpu_custom_instruction_master_start_cpu_fpoint_s1 <= internal_cpu_fpoint_s1_select AND cpu_custom_instruction_master_multi_start;
  --cpu_custom_instruction_master_multi_result mux, which is an e_mux
  cpu_custom_instruction_master_multi_result <= A_REP(internal_cpu_fpoint_s1_select, 32) AND cpu_fpoint_s1_result_from_sa;
  --multi_done mux, which is an e_mux
  cpu_custom_instruction_master_multi_done <= internal_cpu_fpoint_s1_select AND cpu_fpoint_s1_done_from_sa;
  --cpu_custom_instruction_master_reset_n local reset_n, which is an e_assign
  cpu_custom_instruction_master_reset_n <= reset_n;
  --vhdl renameroo for output signals
  cpu_fpoint_s1_select <= internal_cpu_fpoint_s1_select;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpu_data_master_arbitrator is 
        port (
              -- inputs:
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa : IN STD_LOGIC;
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa : IN STD_LOGIC;
                 signal analyzer_input_left_avalon_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                 signal analyzer_input_right_avalon_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                 signal audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal character_buffer_avalon_char_buffer_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal character_buffer_avalon_char_buffer_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal character_buffer_avalon_char_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_byteenable_sdram_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_byteenable_sram_avalon_sram_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                 signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                 signal cpu_data_master_granted_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_data_master_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_compressor_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_compressor_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_compressor_treshold_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_delay_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_delay_decay_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_delay_length_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_master_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_octaver_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_output_power_left_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_output_power_right_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_overdrive_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_overdrive_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_overdrive_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_ps2_avalon_ps2_slave : IN STD_LOGIC;
                 signal cpu_data_master_granted_sdram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_compressor_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_compressor_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_compressor_treshold_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_delay_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_delay_decay_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_delay_length_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_master_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_octaver_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_output_power_left_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_output_power_right_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_ps2_avalon_ps2_slave : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_compressor_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_compressor_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_compressor_treshold_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_delay_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_delay_decay_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_delay_length_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_master_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_octaver_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_output_power_left_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_output_power_right_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                 signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                 signal cpu_data_master_requests_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_data_master_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_compressor_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_compressor_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_compressor_treshold_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_delay_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_delay_decay_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_delay_length_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_master_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_octaver_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_output_power_left_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_output_power_right_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_gain_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_tone_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_volume_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_ps2_avalon_ps2_slave : IN STD_LOGIC;
                 signal cpu_data_master_requests_sdram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer : IN STD_LOGIC;
                 signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer : IN STD_LOGIC;
                 signal d1_analyzer_input_left_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal d1_analyzer_input_right_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer : IN STD_LOGIC;
                 signal d1_character_buffer_avalon_char_buffer_slave_end_xfer : IN STD_LOGIC;
                 signal d1_character_buffer_avalon_char_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal d1_pio_bitcrusher_bypass_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_bitcrusher_crush_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_bitcrusher_downsample_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_bitcrusher_drywet_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_bitcrusher_flavor_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_bitcrusher_tone_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_compressor_bypass_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_compressor_gain_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_compressor_treshold_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_delay_bypass_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_delay_decay_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_delay_length_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_master_volume_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_octaver_bypass_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_octaver_dry_wet_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_output_power_left_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_output_power_right_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_overdrive_asymmetric_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_overdrive_bypass_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_overdrive_gain_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_overdrive_tone_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_overdrive_volume_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_tremolo_stereo_bypass_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_tremolo_stereo_depth_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_tremolo_stereo_mode_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_tremolo_stereo_sweep_a_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pio_tremolo_stereo_sweep_b_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer : IN STD_LOGIC;
                 signal d1_ps2_avalon_ps2_slave_end_xfer : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sram_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal pio_bitcrusher_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_bitcrusher_crush_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pio_bitcrusher_downsample_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pio_bitcrusher_drywet_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_bitcrusher_flavor_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pio_bitcrusher_tone_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_compressor_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_compressor_gain_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pio_compressor_treshold_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_delay_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_delay_decay_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pio_delay_length_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_master_volume_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_octaver_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_octaver_dry_wet_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_output_power_left_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_output_power_right_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_overdrive_asymmetric_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_overdrive_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_overdrive_gain_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_overdrive_tone_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_overdrive_volume_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_tremolo_stereo_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_tremolo_stereo_depth_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_tremolo_stereo_mode_s1_readdata_from_sa : IN STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_a_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pio_tremolo_stereo_sweep_b_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ps2_avalon_ps2_slave_irq_from_sa : IN STD_LOGIC;
                 signal ps2_avalon_ps2_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ps2_avalon_ps2_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : IN STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal sram_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_data_master_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_no_byte_enables_and_last_term : OUT STD_LOGIC;
                 signal cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_data_master_arbitrator;


architecture europa of cpu_data_master_arbitrator is
                signal analyzer_input_left_avalon_slave_readdata_from_sa_part_selected_by_negative_dbs :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal analyzer_input_right_avalon_slave_readdata_from_sa_part_selected_by_negative_dbs :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_data_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_run :  STD_LOGIC;
                signal dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal internal_cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal internal_cpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_data_master_no_byte_enables_and_last_term :  STD_LOGIC;
                signal internal_cpu_data_master_waitrequest :  STD_LOGIC;
                signal last_dbs_term_and_run :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_dbs_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_registered_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal r_3 :  STD_LOGIC;
                signal r_4 :  STD_LOGIC;
                signal r_5 :  STD_LOGIC;
                signal r_6 :  STD_LOGIC;
                signal r_7 :  STD_LOGIC;
                signal registered_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data OR NOT cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control OR NOT cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_analyzer_input_left_avalon_slave OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_analyzer_input_left_avalon_slave OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_analyzer_input_right_avalon_slave OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_analyzer_input_right_avalon_slave OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave OR registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave) OR NOT cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave OR NOT cpu_data_master_read) OR ((registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave AND cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave OR (((registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave AND internal_cpu_data_master_dbs_address(1)) AND internal_cpu_data_master_dbs_address(0)))) OR ((((cpu_data_master_write AND NOT(cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave)) AND internal_cpu_data_master_dbs_address(1)) AND internal_cpu_data_master_dbs_address(0)))) OR NOT cpu_data_master_requests_character_buffer_avalon_char_buffer_slave)))))));
  --cascaded wait assignment, which is an e_assign
  cpu_data_master_run <= ((((((r_0 AND r_1) AND r_2) AND r_3) AND r_4) AND r_5) AND r_6) AND r_7;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave OR NOT cpu_data_master_read) OR (((registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave AND ((internal_cpu_data_master_dbs_address(1) AND internal_cpu_data_master_dbs_address(0)))) AND cpu_data_master_read))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave OR NOT cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT character_buffer_avalon_char_buffer_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_cpu_data_master_dbs_address(1) AND internal_cpu_data_master_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave OR registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave) OR NOT cpu_data_master_requests_character_buffer_avalon_char_control_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave OR NOT cpu_data_master_read) OR ((registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave AND cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_cpu_jtag_debug_module OR NOT cpu_data_master_requests_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_granted_cpu_jtag_debug_module OR NOT cpu_data_master_qualified_request_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_cpu_jtag_debug_module OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_cpu_jtag_debug_module OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave OR NOT cpu_data_master_requests_jtag_uart_avalon_jtag_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 OR NOT cpu_data_master_requests_pio_bitcrusher_bypass_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 OR NOT cpu_data_master_requests_pio_bitcrusher_crush_s1))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 OR NOT cpu_data_master_requests_pio_bitcrusher_downsample_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 OR NOT cpu_data_master_requests_pio_bitcrusher_drywet_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 OR NOT cpu_data_master_requests_pio_bitcrusher_flavor_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 OR NOT cpu_data_master_requests_pio_bitcrusher_tone_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")));
  --r_3 master_run cascaded wait assignment, which is an e_assign
  r_3 <= Vector_To_Std_Logic(((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_compressor_bypass_s1 OR NOT cpu_data_master_requests_pio_compressor_bypass_s1))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_compressor_bypass_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_compressor_bypass_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_compressor_gain_s1 OR NOT cpu_data_master_requests_pio_compressor_gain_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_compressor_gain_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_compressor_gain_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_compressor_treshold_s1 OR NOT cpu_data_master_requests_pio_compressor_treshold_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_compressor_treshold_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_compressor_treshold_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_delay_bypass_s1 OR NOT cpu_data_master_requests_pio_delay_bypass_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_delay_bypass_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_delay_bypass_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_delay_decay_s1 OR NOT cpu_data_master_requests_pio_delay_decay_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_delay_decay_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_delay_decay_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")));
  --r_4 master_run cascaded wait assignment, which is an e_assign
  r_4 <= Vector_To_Std_Logic(((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_delay_length_s1 OR NOT cpu_data_master_requests_pio_delay_length_s1))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_delay_length_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_delay_length_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_master_volume_s1 OR NOT cpu_data_master_requests_pio_master_volume_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_master_volume_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_master_volume_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_octaver_bypass_s1 OR NOT cpu_data_master_requests_pio_octaver_bypass_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_octaver_bypass_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_octaver_bypass_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 OR NOT cpu_data_master_requests_pio_octaver_dry_wet_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_output_power_left_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_output_power_left_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_output_power_right_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))));
  --r_5 master_run cascaded wait assignment, which is an e_assign
  r_5 <= Vector_To_Std_Logic(((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_output_power_right_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 OR NOT cpu_data_master_requests_pio_overdrive_asymmetric_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_overdrive_bypass_s1 OR NOT cpu_data_master_requests_pio_overdrive_bypass_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_bypass_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_bypass_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_overdrive_gain_s1 OR NOT cpu_data_master_requests_pio_overdrive_gain_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_gain_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_gain_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_overdrive_tone_s1 OR NOT cpu_data_master_requests_pio_overdrive_tone_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_tone_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_tone_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_overdrive_volume_s1 OR NOT cpu_data_master_requests_pio_overdrive_volume_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_volume_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))));
  --r_6 master_run cascaded wait assignment, which is an e_assign
  r_6 <= Vector_To_Std_Logic(((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_overdrive_volume_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 OR NOT cpu_data_master_requests_pio_tremolo_stereo_bypass_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 OR NOT cpu_data_master_requests_pio_tremolo_stereo_depth_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 OR NOT cpu_data_master_requests_pio_tremolo_stereo_mode_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 OR NOT cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 OR NOT cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 OR NOT cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read)))))))));
  --r_7 master_run cascaded wait assignment, which is an e_assign
  r_7 <= Vector_To_Std_Logic((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 OR NOT cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave OR registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave) OR NOT cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave OR NOT cpu_data_master_read) OR ((registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave AND cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_data_master_qualified_request_ps2_avalon_ps2_slave OR registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave) OR NOT cpu_data_master_requests_ps2_avalon_ps2_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_data_master_qualified_request_ps2_avalon_ps2_slave OR NOT cpu_data_master_read) OR ((registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave AND cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_ps2_avalon_ps2_slave OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT ps2_avalon_ps2_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((cpu_data_master_qualified_request_sdram_s1 OR ((cpu_data_master_read_data_valid_sdram_s1 AND internal_cpu_data_master_dbs_address(1)))) OR (((cpu_data_master_write AND NOT(or_reduce(cpu_data_master_byteenable_sdram_s1))) AND internal_cpu_data_master_dbs_address(1)))) OR NOT cpu_data_master_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_granted_sdram_s1 OR NOT cpu_data_master_qualified_request_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_data_master_qualified_request_sdram_s1 OR NOT cpu_data_master_read) OR (((cpu_data_master_read_data_valid_sdram_s1 AND (internal_cpu_data_master_dbs_address(1))) AND cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_sdram_s1 OR NOT cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((cpu_data_master_qualified_request_sram_avalon_sram_slave OR ((registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave AND internal_cpu_data_master_dbs_address(1)))) OR (((cpu_data_master_write AND NOT(or_reduce(cpu_data_master_byteenable_sram_avalon_sram_slave))) AND internal_cpu_data_master_dbs_address(1)))) OR NOT cpu_data_master_requests_sram_avalon_sram_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_granted_sram_avalon_sram_slave OR NOT cpu_data_master_qualified_request_sram_avalon_sram_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_data_master_qualified_request_sram_avalon_sram_slave OR NOT cpu_data_master_read) OR (((registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave AND (internal_cpu_data_master_dbs_address(1))) AND cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_sram_avalon_sram_slave OR NOT cpu_data_master_write)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_write)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_data_master_address_to_slave <= cpu_data_master_address(23 DOWNTO 0);
  --unpredictable registered wait state incoming data, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      registered_cpu_data_master_readdata <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      registered_cpu_data_master_readdata <= p1_registered_cpu_data_master_readdata;
    end if;

  end process;

  --registered readdata mux, which is an e_mux
  p1_registered_cpu_data_master_readdata <= ((((A_REP(NOT cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data, 32) OR Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa)) AND ((A_REP(NOT cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control, 32) OR Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_requests_jtag_uart_avalon_jtag_slave, 32) OR jtag_uart_avalon_jtag_slave_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_requests_sdram_s1, 32) OR Std_Logic_Vector'(sdram_s1_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0)));
  --cpu/data_master readdata mux, which is an e_mux
  cpu_data_master_readdata <= ((((((((((((((((((((((((((((((((((((((((A_REP(NOT cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data, 32) OR registered_cpu_data_master_readdata)) AND ((A_REP(NOT cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control, 32) OR registered_cpu_data_master_readdata))) AND ((A_REP(NOT cpu_data_master_requests_analyzer_input_left_avalon_slave, 32) OR analyzer_input_left_avalon_slave_readdata_from_sa_part_selected_by_negative_dbs))) AND ((A_REP(NOT cpu_data_master_requests_analyzer_input_right_avalon_slave, 32) OR analyzer_input_right_avalon_slave_readdata_from_sa_part_selected_by_negative_dbs))) AND ((A_REP(NOT cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave, 32) OR audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_requests_character_buffer_avalon_char_buffer_slave, 32) OR Std_Logic_Vector'(character_buffer_avalon_char_buffer_slave_readdata_from_sa(7 DOWNTO 0) & dbs_8_reg_segment_2 & dbs_8_reg_segment_1 & dbs_8_reg_segment_0)))) AND ((A_REP(NOT cpu_data_master_requests_character_buffer_avalon_char_control_slave, 32) OR character_buffer_avalon_char_control_slave_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_requests_cpu_jtag_debug_module, 32) OR cpu_jtag_debug_module_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_requests_jtag_uart_avalon_jtag_slave, 32) OR registered_cpu_data_master_readdata))) AND ((A_REP(NOT cpu_data_master_requests_pio_bitcrusher_bypass_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_bitcrusher_bypass_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_bitcrusher_crush_s1, 32) OR (std_logic_vector'("0000000000000000000000000000") & (pio_bitcrusher_crush_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_bitcrusher_downsample_s1, 32) OR (std_logic_vector'("000000000000000000000000") & (pio_bitcrusher_downsample_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_bitcrusher_drywet_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_bitcrusher_drywet_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_bitcrusher_flavor_s1, 32) OR (std_logic_vector'("0000000000000000000000000000") & (pio_bitcrusher_flavor_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_bitcrusher_tone_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_bitcrusher_tone_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_compressor_bypass_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_compressor_bypass_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_compressor_gain_s1, 32) OR (std_logic_vector'("000000000000000000000000") & (pio_compressor_gain_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_compressor_treshold_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_compressor_treshold_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_delay_bypass_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_delay_bypass_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_delay_decay_s1, 32) OR (std_logic_vector'("000000000000000000000000") & (pio_delay_decay_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_delay_length_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_delay_length_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_master_volume_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_master_volume_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_octaver_bypass_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_octaver_bypass_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_octaver_dry_wet_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_octaver_dry_wet_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_output_power_left_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_output_power_left_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_output_power_right_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_output_power_right_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_overdrive_asymmetric_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_overdrive_asymmetric_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_overdrive_bypass_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_overdrive_bypass_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_overdrive_gain_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_overdrive_gain_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_overdrive_tone_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_overdrive_tone_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_overdrive_volume_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_overdrive_volume_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_tremolo_stereo_bypass_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_tremolo_stereo_bypass_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_tremolo_stereo_depth_s1, 32) OR (std_logic_vector'("0000000000000000") & (pio_tremolo_stereo_depth_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_tremolo_stereo_mode_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_tremolo_stereo_mode_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1, 32) OR (std_logic_vector'("0000000000000000000000000000") & (pio_tremolo_stereo_sweep_a_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1, 32) OR (std_logic_vector'("0000000000000000000000000000") & (pio_tremolo_stereo_sweep_b_s1_readdata_from_sa))))) AND ((A_REP(NOT cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave, 32) OR pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_requests_ps2_avalon_ps2_slave, 32) OR ps2_avalon_ps2_slave_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_requests_sdram_s1, 32) OR registered_cpu_data_master_readdata))) AND ((A_REP(NOT cpu_data_master_requests_sram_avalon_sram_slave, 32) OR Std_Logic_Vector'(sram_avalon_sram_slave_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0)));
  --actual waitrequest port, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_data_master_waitrequest <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      internal_cpu_data_master_waitrequest <= Vector_To_Std_Logic(NOT (A_WE_StdLogicVector((std_logic'((NOT ((cpu_data_master_read OR cpu_data_master_write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_run AND internal_cpu_data_master_waitrequest))))))));
    end if;

  end process;

  --Negative Dynamic Bus-sizing mux.
  --this mux selects the correct fourth of the 
  --wide data coming from the slave analyzer_input_left/avalon_slave 
  analyzer_input_left_avalon_slave_readdata_from_sa_part_selected_by_negative_dbs <= A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_address_to_slave(3 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000000"))), analyzer_input_left_avalon_slave_readdata_from_sa(31 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_address_to_slave(3 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000001"))), analyzer_input_left_avalon_slave_readdata_from_sa(63 DOWNTO 32), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_address_to_slave(3 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000010"))), analyzer_input_left_avalon_slave_readdata_from_sa(95 DOWNTO 64), analyzer_input_left_avalon_slave_readdata_from_sa(127 DOWNTO 96))));
  --Negative Dynamic Bus-sizing mux.
  --this mux selects the correct fourth of the 
  --wide data coming from the slave analyzer_input_right/avalon_slave 
  analyzer_input_right_avalon_slave_readdata_from_sa_part_selected_by_negative_dbs <= A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_address_to_slave(3 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000000"))), analyzer_input_right_avalon_slave_readdata_from_sa(31 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_address_to_slave(3 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000001"))), analyzer_input_right_avalon_slave_readdata_from_sa(63 DOWNTO 32), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_address_to_slave(3 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000010"))), analyzer_input_right_avalon_slave_readdata_from_sa(95 DOWNTO 64), analyzer_input_right_avalon_slave_readdata_from_sa(127 DOWNTO 96))));
  --no_byte_enables_and_last_term, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_data_master_no_byte_enables_and_last_term <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_cpu_data_master_no_byte_enables_and_last_term <= last_dbs_term_and_run;
    end if;

  end process;

  --compute the last dbs term, which is an e_mux
  last_dbs_term_and_run <= A_WE_StdLogic((std_logic'((cpu_data_master_requests_character_buffer_avalon_char_buffer_slave)) = '1'), (((to_std_logic(((internal_cpu_data_master_dbs_address = std_logic_vector'("11")))) AND cpu_data_master_write) AND NOT(cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave))), A_WE_StdLogic((std_logic'((cpu_data_master_requests_sdram_s1)) = '1'), (((to_std_logic(((internal_cpu_data_master_dbs_address = std_logic_vector'("10")))) AND cpu_data_master_write) AND NOT(or_reduce(cpu_data_master_byteenable_sdram_s1)))), (((to_std_logic(((internal_cpu_data_master_dbs_address = std_logic_vector'("10")))) AND cpu_data_master_write) AND NOT(or_reduce(cpu_data_master_byteenable_sram_avalon_sram_slave))))));
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((((NOT internal_cpu_data_master_no_byte_enables_and_last_term) AND cpu_data_master_requests_character_buffer_avalon_char_buffer_slave) AND cpu_data_master_write) AND NOT(cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave))) OR cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave)))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_character_buffer_avalon_char_buffer_slave AND cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT character_buffer_avalon_char_buffer_slave_waitrequest_from_sa)))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_cpu_data_master_no_byte_enables_and_last_term) AND cpu_data_master_requests_sdram_s1) AND cpu_data_master_write) AND NOT(or_reduce(cpu_data_master_byteenable_sdram_s1)))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read_data_valid_sdram_s1)))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_sdram_s1 AND cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_cpu_data_master_no_byte_enables_and_last_term) AND cpu_data_master_requests_sram_avalon_sram_slave) AND cpu_data_master_write) AND NOT(or_reduce(cpu_data_master_byteenable_sram_avalon_sram_slave)))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_read_data_valid_sram_avalon_sram_slave)))) OR ((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_data_master_granted_sram_avalon_sram_slave AND cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")))));
  --input to dbs-8 stored 0, which is an e_mux
  p1_dbs_8_reg_segment_0 <= character_buffer_avalon_char_buffer_slave_readdata_from_sa;
  --dbs register for dbs-8 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_8_reg_segment_0 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((internal_cpu_data_master_dbs_address(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_8_reg_segment_0 <= p1_dbs_8_reg_segment_0;
      end if;
    end if;

  end process;

  --input to dbs-8 stored 1, which is an e_mux
  p1_dbs_8_reg_segment_1 <= character_buffer_avalon_char_buffer_slave_readdata_from_sa;
  --dbs register for dbs-8 segment 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_8_reg_segment_1 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((internal_cpu_data_master_dbs_address(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000001")))))) = '1' then 
        dbs_8_reg_segment_1 <= p1_dbs_8_reg_segment_1;
      end if;
    end if;

  end process;

  --input to dbs-8 stored 2, which is an e_mux
  p1_dbs_8_reg_segment_2 <= character_buffer_avalon_char_buffer_slave_readdata_from_sa;
  --dbs register for dbs-8 segment 2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_8_reg_segment_2 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((internal_cpu_data_master_dbs_address(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000010")))))) = '1' then 
        dbs_8_reg_segment_2 <= p1_dbs_8_reg_segment_2;
      end if;
    end if;

  end process;

  --mux write dbs 2, which is an e_mux
  cpu_data_master_dbs_write_8 <= A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_writedata(7 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), cpu_data_master_writedata(15 DOWNTO 8), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), cpu_data_master_writedata(23 DOWNTO 16), cpu_data_master_writedata(31 DOWNTO 24))));
  --dbs count increment, which is an e_mux
  cpu_data_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_data_master_requests_character_buffer_avalon_char_buffer_slave)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((cpu_data_master_requests_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((cpu_data_master_requests_sram_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")))), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_cpu_data_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_cpu_data_master_dbs_address)) + (std_logic_vector'("0") & (cpu_data_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= ((pre_dbs_count_enable AND (NOT (((cpu_data_master_requests_character_buffer_avalon_char_buffer_slave AND NOT internal_cpu_data_master_waitrequest) AND cpu_data_master_write)))) AND (NOT ((cpu_data_master_requests_sdram_s1 AND NOT internal_cpu_data_master_waitrequest)))) AND (NOT (((cpu_data_master_requests_sram_avalon_sram_slave AND NOT internal_cpu_data_master_waitrequest) AND cpu_data_master_write)));
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_data_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_cpu_data_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --irq assign, which is an e_assign
  cpu_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(ps2_avalon_ps2_slave_irq_from_sa) & A_ToStdLogicVector(jtag_uart_avalon_jtag_slave_irq_from_sa));
  --input to dbs-16 stored 0, which is an e_mux
  p1_dbs_16_reg_segment_0 <= A_WE_StdLogicVector((std_logic'((cpu_data_master_requests_sdram_s1)) = '1'), sdram_s1_readdata_from_sa, sram_avalon_sram_slave_readdata_from_sa);
  --dbs register for dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_data_master_dbs_address(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
      end if;
    end if;

  end process;

  --mux write dbs 1, which is an e_mux
  cpu_data_master_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_dbs_address(1))) = '1'), cpu_data_master_writedata(31 DOWNTO 16), A_WE_StdLogicVector((std_logic'((NOT (internal_cpu_data_master_dbs_address(1)))) = '1'), cpu_data_master_writedata(15 DOWNTO 0), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_dbs_address(1))) = '1'), cpu_data_master_writedata(31 DOWNTO 16), cpu_data_master_writedata(15 DOWNTO 0))));
  --vhdl renameroo for output signals
  cpu_data_master_address_to_slave <= internal_cpu_data_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_data_master_dbs_address <= internal_cpu_data_master_dbs_address;
  --vhdl renameroo for output signals
  cpu_data_master_no_byte_enables_and_last_term <= internal_cpu_data_master_no_byte_enables_and_last_term;
  --vhdl renameroo for output signals
  cpu_data_master_waitrequest <= internal_cpu_data_master_waitrequest;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_instruction_master_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_instruction_master_granted_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_sram_avalon_sram_slave : IN STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_sram_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sram_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal cpu_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_instruction_master_arbitrator;


architecture europa of cpu_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_instruction_master_address_last_time :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_instruction_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal cpu_instruction_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_instruction_master_read_last_time :  STD_LOGIC;
                signal cpu_instruction_master_run :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal internal_cpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_7 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_cpu_jtag_debug_module OR NOT cpu_instruction_master_requests_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_granted_cpu_jtag_debug_module OR NOT cpu_instruction_master_qualified_request_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_cpu_jtag_debug_module OR NOT cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_instruction_master_run <= r_1 AND r_7;
  --r_7 master_run cascaded wait assignment, which is an e_assign
  r_7 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_sram_avalon_sram_slave OR NOT cpu_instruction_master_requests_sram_avalon_sram_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_granted_sram_avalon_sram_slave OR NOT cpu_instruction_master_qualified_request_sram_avalon_sram_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_sram_avalon_sram_slave OR NOT cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_cpu_instruction_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_read)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_instruction_master_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("110") & cpu_instruction_master_address(20 DOWNTO 0));
  --cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_instruction_master_read_but_no_slave_selected <= (cpu_instruction_master_read AND cpu_instruction_master_run) AND NOT cpu_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_instruction_master_is_granted_some_slave <= cpu_instruction_master_granted_cpu_jtag_debug_module OR cpu_instruction_master_granted_sram_avalon_sram_slave;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_instruction_master_readdatavalid <= cpu_instruction_master_read_data_valid_sram_avalon_sram_slave AND dbs_rdv_counter_overflow;
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_instruction_master_readdatavalid <= (((cpu_instruction_master_read_but_no_slave_selected OR pre_flush_cpu_instruction_master_readdatavalid) OR cpu_instruction_master_read_data_valid_cpu_jtag_debug_module) OR cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_instruction_master_readdatavalid;
  --cpu/instruction_master readdata mux, which is an e_mux
  cpu_instruction_master_readdata <= ((A_REP(NOT ((cpu_instruction_master_qualified_request_cpu_jtag_debug_module AND cpu_instruction_master_read)) , 32) OR cpu_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT cpu_instruction_master_read_data_valid_sram_avalon_sram_slave, 32) OR Std_Logic_Vector'(sram_avalon_sram_slave_readdata_from_sa(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)));
  --actual waitrequest port, which is an e_assign
  internal_cpu_instruction_master_waitrequest <= NOT cpu_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_instruction_master_latency_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      internal_cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_instruction_master_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((cpu_instruction_master_run AND cpu_instruction_master_read))) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_cpu_instruction_master_latency_counter)) /= std_logic_vector'("00")), ((std_logic_vector'("0000000000000000000000000000000") & (internal_cpu_instruction_master_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (A_REP(cpu_instruction_master_requests_sram_avalon_sram_slave, 2))) AND std_logic_vector'("00000000000000000000000000000010")), 2);
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= sram_avalon_sram_slave_readdata_from_sa;
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --dbs count increment, which is an e_mux
  cpu_instruction_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((cpu_instruction_master_requests_sram_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_cpu_instruction_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_cpu_instruction_master_dbs_address)) + (std_logic_vector'("0") & (cpu_instruction_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_instruction_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_cpu_instruction_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  cpu_instruction_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (cpu_instruction_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (cpu_instruction_master_dbs_rdv_counter_inc))), 2);
  --cpu_instruction_master_rdv_inc_mux, which is an e_mux
  cpu_instruction_master_dbs_rdv_counter_inc <= std_logic_vector'("10");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= cpu_instruction_master_read_data_valid_sram_avalon_sram_slave;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_instruction_master_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        cpu_instruction_master_dbs_rdv_counter <= cpu_instruction_master_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= cpu_instruction_master_dbs_rdv_counter(1) AND NOT cpu_instruction_master_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_granted_sram_avalon_sram_slave AND cpu_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")));
  --vhdl renameroo for output signals
  cpu_instruction_master_address_to_slave <= internal_cpu_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_instruction_master_dbs_address <= internal_cpu_instruction_master_dbs_address;
  --vhdl renameroo for output signals
  cpu_instruction_master_latency_counter <= internal_cpu_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  cpu_instruction_master_waitrequest <= internal_cpu_instruction_master_waitrequest;
--synthesis translate_off
    --cpu_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_instruction_master_address_last_time <= std_logic_vector'("000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
      end if;

    end process;

    --cpu/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_instruction_master_waitrequest AND (cpu_instruction_master_read);
      end if;

    end process;

    --cpu_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_instruction_master_address /= cpu_instruction_master_address_last_time))))) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("cpu_instruction_master_address did not heed wait!!!"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
      end if;

    end process;

    --cpu_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_instruction_master_read) /= std_logic'(cpu_instruction_master_read_last_time)))))) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("cpu_instruction_master_read did not heed wait!!!"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpu_fpoint_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                 signal cpu_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal cpu_custom_instruction_master_start_cpu_fpoint_s1 : IN STD_LOGIC;
                 signal cpu_fpoint_s1_done : IN STD_LOGIC;
                 signal cpu_fpoint_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_fpoint_s1_select : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_fpoint_s1_clk_en : OUT STD_LOGIC;
                 signal cpu_fpoint_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_fpoint_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_fpoint_s1_done_from_sa : OUT STD_LOGIC;
                 signal cpu_fpoint_s1_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_fpoint_s1_reset : OUT STD_LOGIC;
                 signal cpu_fpoint_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_fpoint_s1_start : OUT STD_LOGIC
              );
end entity cpu_fpoint_s1_arbitrator;


architecture europa of cpu_fpoint_s1_arbitrator is

begin

  cpu_fpoint_s1_clk_en <= cpu_custom_instruction_master_multi_clk_en;
  cpu_fpoint_s1_dataa <= cpu_custom_instruction_master_multi_dataa;
  cpu_fpoint_s1_datab <= cpu_custom_instruction_master_multi_datab;
  cpu_fpoint_s1_n <= cpu_custom_instruction_master_multi_n (1 DOWNTO 0);
  cpu_fpoint_s1_start <= cpu_custom_instruction_master_start_cpu_fpoint_s1;
  --assign cpu_fpoint_s1_result_from_sa = cpu_fpoint_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_fpoint_s1_result_from_sa <= cpu_fpoint_s1_result;
  --assign cpu_fpoint_s1_done_from_sa = cpu_fpoint_s1_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_fpoint_s1_done_from_sa <= cpu_fpoint_s1_done;
  --cpu_fpoint/s1 local reset_n, which is an e_assign
  cpu_fpoint_s1_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity jtag_uart_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_avalon_jtag_slave_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_jtag_uart_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave);
  --assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readdata_from_sa <= jtag_uart_avalon_jtag_slave_readdata;
  internal_cpu_data_master_requests_jtag_uart_avalon_jtag_slave <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("110100000011000111101000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_avalon_jtag_slave_waitrequest;
  --jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_avalon_jtag_slave_arb_share_set_values <= std_logic_vector'("001");
  --jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (jtag_uart_avalon_jtag_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (jtag_uart_avalon_jtag_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_avalon_jtag_slave_allgrants <= jtag_uart_avalon_jtag_slave_grant_vector;
  --jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_avalon_jtag_slave_waits_for_read OR jtag_uart_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave <= jtag_uart_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND jtag_uart_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 <= or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter_next_value);
  --cpu/data_master jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave <= internal_cpu_data_master_requests_jtag_uart_avalon_jtag_slave AND NOT ((((cpu_data_master_read AND (NOT cpu_data_master_waitrequest))) OR (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write))));
  --jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave <= internal_cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  --cpu/data_master saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  cpu_data_master_saved_grant_jtag_uart_avalon_jtag_slave <= internal_cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  jtag_uart_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_avalon_jtag_slave_chipselect <= internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_read_n <= NOT ((internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave AND cpu_data_master_read));
  --~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_write_n <= NOT ((internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave AND cpu_data_master_write));
  shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_read <= jtag_uart_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_read_cycle <= internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_write <= jtag_uart_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_write_cycle <= internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_irq_from_sa <= jtag_uart_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  cpu_data_master_granted_jtag_uart_avalon_jtag_slave <= internal_cpu_data_master_granted_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave <= internal_cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_jtag_uart_avalon_jtag_slave <= internal_cpu_data_master_requests_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
--synthesis translate_off
    --jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity membuffer_0_avalon_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal membuffer_0_avalon_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal membuffer_0_avalon_master_read : IN STD_LOGIC;
                 signal membuffer_0_avalon_master_write : IN STD_LOGIC;
                 signal membuffer_0_avalon_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal membuffer_0_byteenable_sdram_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal membuffer_0_granted_sdram_s1 : IN STD_LOGIC;
                 signal membuffer_0_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal membuffer_0_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal membuffer_0_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal membuffer_0_requests_sdram_s1 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal membuffer_0_avalon_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal membuffer_0_avalon_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal membuffer_0_avalon_master_reset_n : OUT STD_LOGIC;
                 signal membuffer_0_avalon_master_waitrequest : OUT STD_LOGIC;
                 signal membuffer_0_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal membuffer_0_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity membuffer_0_avalon_master_arbitrator;


architecture europa of membuffer_0_avalon_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal internal_membuffer_0_avalon_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_membuffer_0_avalon_master_waitrequest :  STD_LOGIC;
                signal internal_membuffer_0_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal membuffer_0_avalon_master_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal membuffer_0_avalon_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal membuffer_0_avalon_master_read_last_time :  STD_LOGIC;
                signal membuffer_0_avalon_master_run :  STD_LOGIC;
                signal membuffer_0_avalon_master_write_last_time :  STD_LOGIC;
                signal membuffer_0_avalon_master_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal r_7 :  STD_LOGIC;

begin

  --r_7 master_run cascaded wait assignment, which is an e_assign
  r_7 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((membuffer_0_qualified_request_sdram_s1 OR ((membuffer_0_read_data_valid_sdram_s1 AND internal_membuffer_0_dbs_address(1)))) OR NOT membuffer_0_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((membuffer_0_granted_sdram_s1 OR NOT membuffer_0_qualified_request_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT membuffer_0_qualified_request_sdram_s1 OR NOT membuffer_0_avalon_master_read) OR (((membuffer_0_read_data_valid_sdram_s1 AND (internal_membuffer_0_dbs_address(1))) AND membuffer_0_avalon_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT membuffer_0_qualified_request_sdram_s1 OR NOT membuffer_0_avalon_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_membuffer_0_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(membuffer_0_avalon_master_write)))))))));
  --cascaded wait assignment, which is an e_assign
  membuffer_0_avalon_master_run <= r_7;
  --optimize select-logic by passing only those address bits which matter.
  internal_membuffer_0_avalon_master_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("000000000") & membuffer_0_avalon_master_address(22 DOWNTO 0));
  --input to dbs-16 stored 0, which is an e_mux
  p1_dbs_16_reg_segment_0 <= sdram_s1_readdata_from_sa;
  --dbs register for dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_membuffer_0_dbs_address(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
      end if;
    end if;

  end process;

  --membuffer_0/avalon_master readdata mux, which is an e_mux
  membuffer_0_avalon_master_readdata <= Std_Logic_Vector'(sdram_s1_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0);
  --mux write dbs 1, which is an e_mux
  membuffer_0_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_membuffer_0_dbs_address(1))) = '1'), membuffer_0_avalon_master_writedata(31 DOWNTO 16), membuffer_0_avalon_master_writedata(15 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_membuffer_0_avalon_master_waitrequest <= NOT membuffer_0_avalon_master_run;
  --membuffer_0_avalon_master_reset_n assignment, which is an e_assign
  membuffer_0_avalon_master_reset_n <= reset_n;
  --dbs count increment, which is an e_mux
  membuffer_0_avalon_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((membuffer_0_requests_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_membuffer_0_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_membuffer_0_dbs_address)) + (std_logic_vector'("0") & (membuffer_0_avalon_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_membuffer_0_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_membuffer_0_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(membuffer_0_read_data_valid_sdram_s1))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((membuffer_0_granted_sdram_s1 AND membuffer_0_avalon_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))))));
  --vhdl renameroo for output signals
  membuffer_0_avalon_master_address_to_slave <= internal_membuffer_0_avalon_master_address_to_slave;
  --vhdl renameroo for output signals
  membuffer_0_avalon_master_waitrequest <= internal_membuffer_0_avalon_master_waitrequest;
  --vhdl renameroo for output signals
  membuffer_0_dbs_address <= internal_membuffer_0_dbs_address;
--synthesis translate_off
    --membuffer_0_avalon_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        membuffer_0_avalon_master_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        membuffer_0_avalon_master_address_last_time <= membuffer_0_avalon_master_address;
      end if;

    end process;

    --membuffer_0/avalon_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_membuffer_0_avalon_master_waitrequest AND ((membuffer_0_avalon_master_read OR membuffer_0_avalon_master_write));
      end if;

    end process;

    --membuffer_0_avalon_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((membuffer_0_avalon_master_address /= membuffer_0_avalon_master_address_last_time))))) = '1' then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("membuffer_0_avalon_master_address did not heed wait!!!"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --membuffer_0_avalon_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        membuffer_0_avalon_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        membuffer_0_avalon_master_read_last_time <= membuffer_0_avalon_master_read;
      end if;

    end process;

    --membuffer_0_avalon_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(membuffer_0_avalon_master_read) /= std_logic'(membuffer_0_avalon_master_read_last_time)))))) = '1' then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("membuffer_0_avalon_master_read did not heed wait!!!"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --membuffer_0_avalon_master_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        membuffer_0_avalon_master_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        membuffer_0_avalon_master_write_last_time <= membuffer_0_avalon_master_write;
      end if;

    end process;

    --membuffer_0_avalon_master_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(membuffer_0_avalon_master_write) /= std_logic'(membuffer_0_avalon_master_write_last_time)))))) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("membuffer_0_avalon_master_write did not heed wait!!!"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --membuffer_0_avalon_master_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        membuffer_0_avalon_master_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        membuffer_0_avalon_master_writedata_last_time <= membuffer_0_avalon_master_writedata;
      end if;

    end process;

    --membuffer_0_avalon_master_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((membuffer_0_avalon_master_writedata /= membuffer_0_avalon_master_writedata_last_time)))) AND membuffer_0_avalon_master_write)) = '1' then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("membuffer_0_avalon_master_writedata did not heed wait!!!"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_bitcrusher_bypass_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_bitcrusher_bypass_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                 signal d1_pio_bitcrusher_bypass_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_bitcrusher_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_bitcrusher_bypass_s1_chipselect : OUT STD_LOGIC;
                 signal pio_bitcrusher_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_bitcrusher_bypass_s1_reset_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_bypass_s1_write_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_bypass_s1_writedata : OUT STD_LOGIC
              );
end entity pio_bitcrusher_bypass_s1_arbitrator;


architecture europa of pio_bitcrusher_bypass_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_allgrants :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_any_continuerequest :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_bypass_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_bypass_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_bypass_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_begins_xfer :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_end_xfer :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_grant_vector :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_waits_for_read :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_bitcrusher_bypass_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_bitcrusher_bypass_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_bitcrusher_bypass_s1_end_xfer;
    end if;

  end process;

  pio_bitcrusher_bypass_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1);
  --assign pio_bitcrusher_bypass_s1_readdata_from_sa = pio_bitcrusher_bypass_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_bitcrusher_bypass_s1_readdata_from_sa <= pio_bitcrusher_bypass_s1_readdata;
  internal_cpu_data_master_requests_pio_bitcrusher_bypass_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000011110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_bitcrusher_bypass_s1_arb_share_counter set values, which is an e_mux
  pio_bitcrusher_bypass_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_bitcrusher_bypass_s1_non_bursting_master_requests mux, which is an e_mux
  pio_bitcrusher_bypass_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_bitcrusher_bypass_s1;
  --pio_bitcrusher_bypass_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_bitcrusher_bypass_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_bitcrusher_bypass_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_bitcrusher_bypass_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_bitcrusher_bypass_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_bypass_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_bitcrusher_bypass_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_bypass_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_bitcrusher_bypass_s1_allgrants all slave grants, which is an e_mux
  pio_bitcrusher_bypass_s1_allgrants <= pio_bitcrusher_bypass_s1_grant_vector;
  --pio_bitcrusher_bypass_s1_end_xfer assignment, which is an e_assign
  pio_bitcrusher_bypass_s1_end_xfer <= NOT ((pio_bitcrusher_bypass_s1_waits_for_read OR pio_bitcrusher_bypass_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_bitcrusher_bypass_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_bitcrusher_bypass_s1 <= pio_bitcrusher_bypass_s1_end_xfer AND (((NOT pio_bitcrusher_bypass_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_bitcrusher_bypass_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_bitcrusher_bypass_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_bitcrusher_bypass_s1 AND pio_bitcrusher_bypass_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_bypass_s1 AND NOT pio_bitcrusher_bypass_s1_non_bursting_master_requests));
  --pio_bitcrusher_bypass_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_bypass_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_bypass_s1_arb_counter_enable) = '1' then 
        pio_bitcrusher_bypass_s1_arb_share_counter <= pio_bitcrusher_bypass_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_bitcrusher_bypass_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_bypass_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_bitcrusher_bypass_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_bitcrusher_bypass_s1)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_bypass_s1 AND NOT pio_bitcrusher_bypass_s1_non_bursting_master_requests)))) = '1' then 
        pio_bitcrusher_bypass_s1_slavearbiterlockenable <= or_reduce(pio_bitcrusher_bypass_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_bitcrusher_bypass/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_bitcrusher_bypass_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_bitcrusher_bypass_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_bitcrusher_bypass_s1_slavearbiterlockenable2 <= or_reduce(pio_bitcrusher_bypass_s1_arb_share_counter_next_value);
  --cpu/data_master pio_bitcrusher_bypass/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_bitcrusher_bypass_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_bitcrusher_bypass_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_bitcrusher_bypass_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_bypass_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_bitcrusher_bypass_s1_writedata mux, which is an e_mux
  pio_bitcrusher_bypass_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_bitcrusher_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1;
  --cpu/data_master saved-grant pio_bitcrusher_bypass/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_bitcrusher_bypass_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_bypass_s1;
  --allow new arb cycle for pio_bitcrusher_bypass/s1, which is an e_assign
  pio_bitcrusher_bypass_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_bitcrusher_bypass_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_bitcrusher_bypass_s1_master_qreq_vector <= std_logic'('1');
  --pio_bitcrusher_bypass_s1_reset_n assignment, which is an e_assign
  pio_bitcrusher_bypass_s1_reset_n <= reset_n;
  pio_bitcrusher_bypass_s1_chipselect <= internal_cpu_data_master_granted_pio_bitcrusher_bypass_s1;
  --pio_bitcrusher_bypass_s1_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_bypass_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_bitcrusher_bypass_s1_begins_xfer) = '1'), pio_bitcrusher_bypass_s1_unreg_firsttransfer, pio_bitcrusher_bypass_s1_reg_firsttransfer);
  --pio_bitcrusher_bypass_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_bypass_s1_unreg_firsttransfer <= NOT ((pio_bitcrusher_bypass_s1_slavearbiterlockenable AND pio_bitcrusher_bypass_s1_any_continuerequest));
  --pio_bitcrusher_bypass_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_bypass_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_bypass_s1_begins_xfer) = '1' then 
        pio_bitcrusher_bypass_s1_reg_firsttransfer <= pio_bitcrusher_bypass_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_bitcrusher_bypass_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_bitcrusher_bypass_s1_beginbursttransfer_internal <= pio_bitcrusher_bypass_s1_begins_xfer;
  --~pio_bitcrusher_bypass_s1_write_n assignment, which is an e_mux
  pio_bitcrusher_bypass_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_bitcrusher_bypass_s1 AND cpu_data_master_write));
  shifted_address_to_pio_bitcrusher_bypass_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_bitcrusher_bypass_s1_address mux, which is an e_mux
  pio_bitcrusher_bypass_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_bitcrusher_bypass_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_bitcrusher_bypass_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_bitcrusher_bypass_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_bitcrusher_bypass_s1_end_xfer <= pio_bitcrusher_bypass_s1_end_xfer;
    end if;

  end process;

  --pio_bitcrusher_bypass_s1_waits_for_read in a cycle, which is an e_mux
  pio_bitcrusher_bypass_s1_waits_for_read <= pio_bitcrusher_bypass_s1_in_a_read_cycle AND pio_bitcrusher_bypass_s1_begins_xfer;
  --pio_bitcrusher_bypass_s1_in_a_read_cycle assignment, which is an e_assign
  pio_bitcrusher_bypass_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_bypass_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_bitcrusher_bypass_s1_in_a_read_cycle;
  --pio_bitcrusher_bypass_s1_waits_for_write in a cycle, which is an e_mux
  pio_bitcrusher_bypass_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_bitcrusher_bypass_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_bitcrusher_bypass_s1_in_a_write_cycle assignment, which is an e_assign
  pio_bitcrusher_bypass_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_bypass_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_bitcrusher_bypass_s1_in_a_write_cycle;
  wait_for_pio_bitcrusher_bypass_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_bitcrusher_bypass_s1 <= internal_cpu_data_master_granted_pio_bitcrusher_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_bitcrusher_bypass_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_bypass_s1;
--synthesis translate_off
    --pio_bitcrusher_bypass/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_bitcrusher_crush_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_bitcrusher_crush_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                 signal d1_pio_bitcrusher_crush_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_bitcrusher_crush_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_bitcrusher_crush_s1_chipselect : OUT STD_LOGIC;
                 signal pio_bitcrusher_crush_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pio_bitcrusher_crush_s1_reset_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_crush_s1_write_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_crush_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
              );
end entity pio_bitcrusher_crush_s1_arbitrator;


architecture europa of pio_bitcrusher_crush_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_allgrants :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_any_continuerequest :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_crush_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_crush_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_crush_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_begins_xfer :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_end_xfer :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_grant_vector :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_waits_for_read :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_bitcrusher_crush_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_bitcrusher_crush_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_bitcrusher_crush_s1_end_xfer;
    end if;

  end process;

  pio_bitcrusher_crush_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_bitcrusher_crush_s1);
  --assign pio_bitcrusher_crush_s1_readdata_from_sa = pio_bitcrusher_crush_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_bitcrusher_crush_s1_readdata_from_sa <= pio_bitcrusher_crush_s1_readdata;
  internal_cpu_data_master_requests_pio_bitcrusher_crush_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000100000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_bitcrusher_crush_s1_arb_share_counter set values, which is an e_mux
  pio_bitcrusher_crush_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_bitcrusher_crush_s1_non_bursting_master_requests mux, which is an e_mux
  pio_bitcrusher_crush_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_bitcrusher_crush_s1;
  --pio_bitcrusher_crush_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_bitcrusher_crush_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_bitcrusher_crush_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_bitcrusher_crush_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_bitcrusher_crush_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_crush_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_bitcrusher_crush_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_crush_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_bitcrusher_crush_s1_allgrants all slave grants, which is an e_mux
  pio_bitcrusher_crush_s1_allgrants <= pio_bitcrusher_crush_s1_grant_vector;
  --pio_bitcrusher_crush_s1_end_xfer assignment, which is an e_assign
  pio_bitcrusher_crush_s1_end_xfer <= NOT ((pio_bitcrusher_crush_s1_waits_for_read OR pio_bitcrusher_crush_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_bitcrusher_crush_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_bitcrusher_crush_s1 <= pio_bitcrusher_crush_s1_end_xfer AND (((NOT pio_bitcrusher_crush_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_bitcrusher_crush_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_bitcrusher_crush_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_bitcrusher_crush_s1 AND pio_bitcrusher_crush_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_crush_s1 AND NOT pio_bitcrusher_crush_s1_non_bursting_master_requests));
  --pio_bitcrusher_crush_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_crush_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_crush_s1_arb_counter_enable) = '1' then 
        pio_bitcrusher_crush_s1_arb_share_counter <= pio_bitcrusher_crush_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_bitcrusher_crush_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_crush_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_bitcrusher_crush_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_bitcrusher_crush_s1)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_crush_s1 AND NOT pio_bitcrusher_crush_s1_non_bursting_master_requests)))) = '1' then 
        pio_bitcrusher_crush_s1_slavearbiterlockenable <= or_reduce(pio_bitcrusher_crush_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_bitcrusher_crush/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_bitcrusher_crush_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_bitcrusher_crush_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_bitcrusher_crush_s1_slavearbiterlockenable2 <= or_reduce(pio_bitcrusher_crush_s1_arb_share_counter_next_value);
  --cpu/data_master pio_bitcrusher_crush/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_bitcrusher_crush_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_bitcrusher_crush_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_bitcrusher_crush_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_crush_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_bitcrusher_crush_s1_writedata mux, which is an e_mux
  pio_bitcrusher_crush_s1_writedata <= cpu_data_master_writedata (3 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_bitcrusher_crush_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_crush_s1;
  --cpu/data_master saved-grant pio_bitcrusher_crush/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_bitcrusher_crush_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_crush_s1;
  --allow new arb cycle for pio_bitcrusher_crush/s1, which is an e_assign
  pio_bitcrusher_crush_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_bitcrusher_crush_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_bitcrusher_crush_s1_master_qreq_vector <= std_logic'('1');
  --pio_bitcrusher_crush_s1_reset_n assignment, which is an e_assign
  pio_bitcrusher_crush_s1_reset_n <= reset_n;
  pio_bitcrusher_crush_s1_chipselect <= internal_cpu_data_master_granted_pio_bitcrusher_crush_s1;
  --pio_bitcrusher_crush_s1_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_crush_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_bitcrusher_crush_s1_begins_xfer) = '1'), pio_bitcrusher_crush_s1_unreg_firsttransfer, pio_bitcrusher_crush_s1_reg_firsttransfer);
  --pio_bitcrusher_crush_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_crush_s1_unreg_firsttransfer <= NOT ((pio_bitcrusher_crush_s1_slavearbiterlockenable AND pio_bitcrusher_crush_s1_any_continuerequest));
  --pio_bitcrusher_crush_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_crush_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_crush_s1_begins_xfer) = '1' then 
        pio_bitcrusher_crush_s1_reg_firsttransfer <= pio_bitcrusher_crush_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_bitcrusher_crush_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_bitcrusher_crush_s1_beginbursttransfer_internal <= pio_bitcrusher_crush_s1_begins_xfer;
  --~pio_bitcrusher_crush_s1_write_n assignment, which is an e_mux
  pio_bitcrusher_crush_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_bitcrusher_crush_s1 AND cpu_data_master_write));
  shifted_address_to_pio_bitcrusher_crush_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_bitcrusher_crush_s1_address mux, which is an e_mux
  pio_bitcrusher_crush_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_bitcrusher_crush_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_bitcrusher_crush_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_bitcrusher_crush_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_bitcrusher_crush_s1_end_xfer <= pio_bitcrusher_crush_s1_end_xfer;
    end if;

  end process;

  --pio_bitcrusher_crush_s1_waits_for_read in a cycle, which is an e_mux
  pio_bitcrusher_crush_s1_waits_for_read <= pio_bitcrusher_crush_s1_in_a_read_cycle AND pio_bitcrusher_crush_s1_begins_xfer;
  --pio_bitcrusher_crush_s1_in_a_read_cycle assignment, which is an e_assign
  pio_bitcrusher_crush_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_crush_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_bitcrusher_crush_s1_in_a_read_cycle;
  --pio_bitcrusher_crush_s1_waits_for_write in a cycle, which is an e_mux
  pio_bitcrusher_crush_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_bitcrusher_crush_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_bitcrusher_crush_s1_in_a_write_cycle assignment, which is an e_assign
  pio_bitcrusher_crush_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_crush_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_bitcrusher_crush_s1_in_a_write_cycle;
  wait_for_pio_bitcrusher_crush_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_bitcrusher_crush_s1 <= internal_cpu_data_master_granted_pio_bitcrusher_crush_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_crush_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_bitcrusher_crush_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_crush_s1;
--synthesis translate_off
    --pio_bitcrusher_crush/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_bitcrusher_downsample_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_bitcrusher_downsample_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                 signal d1_pio_bitcrusher_downsample_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_bitcrusher_downsample_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_bitcrusher_downsample_s1_chipselect : OUT STD_LOGIC;
                 signal pio_bitcrusher_downsample_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pio_bitcrusher_downsample_s1_reset_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_downsample_s1_write_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_downsample_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity pio_bitcrusher_downsample_s1_arbitrator;


architecture europa of pio_bitcrusher_downsample_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_allgrants :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_any_continuerequest :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_downsample_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_downsample_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_downsample_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_begins_xfer :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_end_xfer :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_grant_vector :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_pretend_byte_enable :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_waits_for_read :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_bitcrusher_downsample_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_bitcrusher_downsample_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_bitcrusher_downsample_s1_end_xfer;
    end if;

  end process;

  pio_bitcrusher_downsample_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1);
  --assign pio_bitcrusher_downsample_s1_readdata_from_sa = pio_bitcrusher_downsample_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_bitcrusher_downsample_s1_readdata_from_sa <= pio_bitcrusher_downsample_s1_readdata;
  internal_cpu_data_master_requests_pio_bitcrusher_downsample_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000100010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_bitcrusher_downsample_s1_arb_share_counter set values, which is an e_mux
  pio_bitcrusher_downsample_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_bitcrusher_downsample_s1_non_bursting_master_requests mux, which is an e_mux
  pio_bitcrusher_downsample_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_bitcrusher_downsample_s1;
  --pio_bitcrusher_downsample_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_bitcrusher_downsample_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_bitcrusher_downsample_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_bitcrusher_downsample_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_bitcrusher_downsample_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_downsample_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_bitcrusher_downsample_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_downsample_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_bitcrusher_downsample_s1_allgrants all slave grants, which is an e_mux
  pio_bitcrusher_downsample_s1_allgrants <= pio_bitcrusher_downsample_s1_grant_vector;
  --pio_bitcrusher_downsample_s1_end_xfer assignment, which is an e_assign
  pio_bitcrusher_downsample_s1_end_xfer <= NOT ((pio_bitcrusher_downsample_s1_waits_for_read OR pio_bitcrusher_downsample_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_bitcrusher_downsample_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_bitcrusher_downsample_s1 <= pio_bitcrusher_downsample_s1_end_xfer AND (((NOT pio_bitcrusher_downsample_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_bitcrusher_downsample_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_bitcrusher_downsample_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_bitcrusher_downsample_s1 AND pio_bitcrusher_downsample_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_downsample_s1 AND NOT pio_bitcrusher_downsample_s1_non_bursting_master_requests));
  --pio_bitcrusher_downsample_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_downsample_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_downsample_s1_arb_counter_enable) = '1' then 
        pio_bitcrusher_downsample_s1_arb_share_counter <= pio_bitcrusher_downsample_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_bitcrusher_downsample_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_downsample_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_bitcrusher_downsample_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_bitcrusher_downsample_s1)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_downsample_s1 AND NOT pio_bitcrusher_downsample_s1_non_bursting_master_requests)))) = '1' then 
        pio_bitcrusher_downsample_s1_slavearbiterlockenable <= or_reduce(pio_bitcrusher_downsample_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_bitcrusher_downsample/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_bitcrusher_downsample_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_bitcrusher_downsample_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_bitcrusher_downsample_s1_slavearbiterlockenable2 <= or_reduce(pio_bitcrusher_downsample_s1_arb_share_counter_next_value);
  --cpu/data_master pio_bitcrusher_downsample/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_bitcrusher_downsample_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_bitcrusher_downsample_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_bitcrusher_downsample_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_downsample_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_bitcrusher_downsample_s1_writedata mux, which is an e_mux
  pio_bitcrusher_downsample_s1_writedata <= cpu_data_master_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1;
  --cpu/data_master saved-grant pio_bitcrusher_downsample/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_bitcrusher_downsample_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_downsample_s1;
  --allow new arb cycle for pio_bitcrusher_downsample/s1, which is an e_assign
  pio_bitcrusher_downsample_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_bitcrusher_downsample_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_bitcrusher_downsample_s1_master_qreq_vector <= std_logic'('1');
  --pio_bitcrusher_downsample_s1_reset_n assignment, which is an e_assign
  pio_bitcrusher_downsample_s1_reset_n <= reset_n;
  pio_bitcrusher_downsample_s1_chipselect <= internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1;
  --pio_bitcrusher_downsample_s1_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_downsample_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_bitcrusher_downsample_s1_begins_xfer) = '1'), pio_bitcrusher_downsample_s1_unreg_firsttransfer, pio_bitcrusher_downsample_s1_reg_firsttransfer);
  --pio_bitcrusher_downsample_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_downsample_s1_unreg_firsttransfer <= NOT ((pio_bitcrusher_downsample_s1_slavearbiterlockenable AND pio_bitcrusher_downsample_s1_any_continuerequest));
  --pio_bitcrusher_downsample_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_downsample_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_downsample_s1_begins_xfer) = '1' then 
        pio_bitcrusher_downsample_s1_reg_firsttransfer <= pio_bitcrusher_downsample_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_bitcrusher_downsample_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_bitcrusher_downsample_s1_beginbursttransfer_internal <= pio_bitcrusher_downsample_s1_begins_xfer;
  --~pio_bitcrusher_downsample_s1_write_n assignment, which is an e_mux
  pio_bitcrusher_downsample_s1_write_n <= NOT ((((internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1 AND cpu_data_master_write)) AND pio_bitcrusher_downsample_s1_pretend_byte_enable));
  shifted_address_to_pio_bitcrusher_downsample_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_bitcrusher_downsample_s1_address mux, which is an e_mux
  pio_bitcrusher_downsample_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_bitcrusher_downsample_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_bitcrusher_downsample_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_bitcrusher_downsample_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_bitcrusher_downsample_s1_end_xfer <= pio_bitcrusher_downsample_s1_end_xfer;
    end if;

  end process;

  --pio_bitcrusher_downsample_s1_waits_for_read in a cycle, which is an e_mux
  pio_bitcrusher_downsample_s1_waits_for_read <= pio_bitcrusher_downsample_s1_in_a_read_cycle AND pio_bitcrusher_downsample_s1_begins_xfer;
  --pio_bitcrusher_downsample_s1_in_a_read_cycle assignment, which is an e_assign
  pio_bitcrusher_downsample_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_bitcrusher_downsample_s1_in_a_read_cycle;
  --pio_bitcrusher_downsample_s1_waits_for_write in a cycle, which is an e_mux
  pio_bitcrusher_downsample_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_bitcrusher_downsample_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_bitcrusher_downsample_s1_in_a_write_cycle assignment, which is an e_assign
  pio_bitcrusher_downsample_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_bitcrusher_downsample_s1_in_a_write_cycle;
  wait_for_pio_bitcrusher_downsample_s1_counter <= std_logic'('0');
  --pio_bitcrusher_downsample_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  pio_bitcrusher_downsample_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_bitcrusher_downsample_s1 <= internal_cpu_data_master_granted_pio_bitcrusher_downsample_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_bitcrusher_downsample_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_downsample_s1;
--synthesis translate_off
    --pio_bitcrusher_downsample/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_bitcrusher_drywet_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_bitcrusher_drywet_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                 signal d1_pio_bitcrusher_drywet_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_bitcrusher_drywet_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_bitcrusher_drywet_s1_chipselect : OUT STD_LOGIC;
                 signal pio_bitcrusher_drywet_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_bitcrusher_drywet_s1_reset_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_drywet_s1_write_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_drywet_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_bitcrusher_drywet_s1_arbitrator;


architecture europa of pio_bitcrusher_drywet_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_allgrants :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_any_continuerequest :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_drywet_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_drywet_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_drywet_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_begins_xfer :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_end_xfer :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_grant_vector :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_waits_for_read :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_bitcrusher_drywet_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_bitcrusher_drywet_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_bitcrusher_drywet_s1_end_xfer;
    end if;

  end process;

  pio_bitcrusher_drywet_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1);
  --assign pio_bitcrusher_drywet_s1_readdata_from_sa = pio_bitcrusher_drywet_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_bitcrusher_drywet_s1_readdata_from_sa <= pio_bitcrusher_drywet_s1_readdata;
  internal_cpu_data_master_requests_pio_bitcrusher_drywet_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000100100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_bitcrusher_drywet_s1_arb_share_counter set values, which is an e_mux
  pio_bitcrusher_drywet_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_bitcrusher_drywet_s1_non_bursting_master_requests mux, which is an e_mux
  pio_bitcrusher_drywet_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_bitcrusher_drywet_s1;
  --pio_bitcrusher_drywet_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_bitcrusher_drywet_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_bitcrusher_drywet_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_bitcrusher_drywet_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_bitcrusher_drywet_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_drywet_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_bitcrusher_drywet_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_drywet_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_bitcrusher_drywet_s1_allgrants all slave grants, which is an e_mux
  pio_bitcrusher_drywet_s1_allgrants <= pio_bitcrusher_drywet_s1_grant_vector;
  --pio_bitcrusher_drywet_s1_end_xfer assignment, which is an e_assign
  pio_bitcrusher_drywet_s1_end_xfer <= NOT ((pio_bitcrusher_drywet_s1_waits_for_read OR pio_bitcrusher_drywet_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_bitcrusher_drywet_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_bitcrusher_drywet_s1 <= pio_bitcrusher_drywet_s1_end_xfer AND (((NOT pio_bitcrusher_drywet_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_bitcrusher_drywet_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_bitcrusher_drywet_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_bitcrusher_drywet_s1 AND pio_bitcrusher_drywet_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_drywet_s1 AND NOT pio_bitcrusher_drywet_s1_non_bursting_master_requests));
  --pio_bitcrusher_drywet_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_drywet_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_drywet_s1_arb_counter_enable) = '1' then 
        pio_bitcrusher_drywet_s1_arb_share_counter <= pio_bitcrusher_drywet_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_bitcrusher_drywet_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_drywet_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_bitcrusher_drywet_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_bitcrusher_drywet_s1)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_drywet_s1 AND NOT pio_bitcrusher_drywet_s1_non_bursting_master_requests)))) = '1' then 
        pio_bitcrusher_drywet_s1_slavearbiterlockenable <= or_reduce(pio_bitcrusher_drywet_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_bitcrusher_drywet/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_bitcrusher_drywet_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_bitcrusher_drywet_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_bitcrusher_drywet_s1_slavearbiterlockenable2 <= or_reduce(pio_bitcrusher_drywet_s1_arb_share_counter_next_value);
  --cpu/data_master pio_bitcrusher_drywet/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_bitcrusher_drywet_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_bitcrusher_drywet_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_bitcrusher_drywet_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_drywet_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_bitcrusher_drywet_s1_writedata mux, which is an e_mux
  pio_bitcrusher_drywet_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_bitcrusher_drywet_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1;
  --cpu/data_master saved-grant pio_bitcrusher_drywet/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_bitcrusher_drywet_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_drywet_s1;
  --allow new arb cycle for pio_bitcrusher_drywet/s1, which is an e_assign
  pio_bitcrusher_drywet_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_bitcrusher_drywet_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_bitcrusher_drywet_s1_master_qreq_vector <= std_logic'('1');
  --pio_bitcrusher_drywet_s1_reset_n assignment, which is an e_assign
  pio_bitcrusher_drywet_s1_reset_n <= reset_n;
  pio_bitcrusher_drywet_s1_chipselect <= internal_cpu_data_master_granted_pio_bitcrusher_drywet_s1;
  --pio_bitcrusher_drywet_s1_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_drywet_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_bitcrusher_drywet_s1_begins_xfer) = '1'), pio_bitcrusher_drywet_s1_unreg_firsttransfer, pio_bitcrusher_drywet_s1_reg_firsttransfer);
  --pio_bitcrusher_drywet_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_drywet_s1_unreg_firsttransfer <= NOT ((pio_bitcrusher_drywet_s1_slavearbiterlockenable AND pio_bitcrusher_drywet_s1_any_continuerequest));
  --pio_bitcrusher_drywet_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_drywet_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_drywet_s1_begins_xfer) = '1' then 
        pio_bitcrusher_drywet_s1_reg_firsttransfer <= pio_bitcrusher_drywet_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_bitcrusher_drywet_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_bitcrusher_drywet_s1_beginbursttransfer_internal <= pio_bitcrusher_drywet_s1_begins_xfer;
  --~pio_bitcrusher_drywet_s1_write_n assignment, which is an e_mux
  pio_bitcrusher_drywet_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_bitcrusher_drywet_s1 AND cpu_data_master_write));
  shifted_address_to_pio_bitcrusher_drywet_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_bitcrusher_drywet_s1_address mux, which is an e_mux
  pio_bitcrusher_drywet_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_bitcrusher_drywet_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_bitcrusher_drywet_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_bitcrusher_drywet_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_bitcrusher_drywet_s1_end_xfer <= pio_bitcrusher_drywet_s1_end_xfer;
    end if;

  end process;

  --pio_bitcrusher_drywet_s1_waits_for_read in a cycle, which is an e_mux
  pio_bitcrusher_drywet_s1_waits_for_read <= pio_bitcrusher_drywet_s1_in_a_read_cycle AND pio_bitcrusher_drywet_s1_begins_xfer;
  --pio_bitcrusher_drywet_s1_in_a_read_cycle assignment, which is an e_assign
  pio_bitcrusher_drywet_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_drywet_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_bitcrusher_drywet_s1_in_a_read_cycle;
  --pio_bitcrusher_drywet_s1_waits_for_write in a cycle, which is an e_mux
  pio_bitcrusher_drywet_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_bitcrusher_drywet_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_bitcrusher_drywet_s1_in_a_write_cycle assignment, which is an e_assign
  pio_bitcrusher_drywet_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_drywet_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_bitcrusher_drywet_s1_in_a_write_cycle;
  wait_for_pio_bitcrusher_drywet_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_bitcrusher_drywet_s1 <= internal_cpu_data_master_granted_pio_bitcrusher_drywet_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_bitcrusher_drywet_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_drywet_s1;
--synthesis translate_off
    --pio_bitcrusher_drywet/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_bitcrusher_flavor_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_bitcrusher_flavor_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                 signal d1_pio_bitcrusher_flavor_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_bitcrusher_flavor_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_bitcrusher_flavor_s1_chipselect : OUT STD_LOGIC;
                 signal pio_bitcrusher_flavor_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pio_bitcrusher_flavor_s1_reset_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_flavor_s1_write_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_flavor_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
              );
end entity pio_bitcrusher_flavor_s1_arbitrator;


architecture europa of pio_bitcrusher_flavor_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_allgrants :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_any_continuerequest :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_flavor_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_flavor_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_flavor_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_begins_xfer :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_end_xfer :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_grant_vector :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_waits_for_read :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_bitcrusher_flavor_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_bitcrusher_flavor_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_bitcrusher_flavor_s1_end_xfer;
    end if;

  end process;

  pio_bitcrusher_flavor_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1);
  --assign pio_bitcrusher_flavor_s1_readdata_from_sa = pio_bitcrusher_flavor_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_bitcrusher_flavor_s1_readdata_from_sa <= pio_bitcrusher_flavor_s1_readdata;
  internal_cpu_data_master_requests_pio_bitcrusher_flavor_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000111010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_bitcrusher_flavor_s1_arb_share_counter set values, which is an e_mux
  pio_bitcrusher_flavor_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_bitcrusher_flavor_s1_non_bursting_master_requests mux, which is an e_mux
  pio_bitcrusher_flavor_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_bitcrusher_flavor_s1;
  --pio_bitcrusher_flavor_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_bitcrusher_flavor_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_bitcrusher_flavor_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_bitcrusher_flavor_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_bitcrusher_flavor_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_flavor_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_bitcrusher_flavor_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_flavor_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_bitcrusher_flavor_s1_allgrants all slave grants, which is an e_mux
  pio_bitcrusher_flavor_s1_allgrants <= pio_bitcrusher_flavor_s1_grant_vector;
  --pio_bitcrusher_flavor_s1_end_xfer assignment, which is an e_assign
  pio_bitcrusher_flavor_s1_end_xfer <= NOT ((pio_bitcrusher_flavor_s1_waits_for_read OR pio_bitcrusher_flavor_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_bitcrusher_flavor_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_bitcrusher_flavor_s1 <= pio_bitcrusher_flavor_s1_end_xfer AND (((NOT pio_bitcrusher_flavor_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_bitcrusher_flavor_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_bitcrusher_flavor_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_bitcrusher_flavor_s1 AND pio_bitcrusher_flavor_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_flavor_s1 AND NOT pio_bitcrusher_flavor_s1_non_bursting_master_requests));
  --pio_bitcrusher_flavor_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_flavor_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_flavor_s1_arb_counter_enable) = '1' then 
        pio_bitcrusher_flavor_s1_arb_share_counter <= pio_bitcrusher_flavor_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_bitcrusher_flavor_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_flavor_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_bitcrusher_flavor_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_bitcrusher_flavor_s1)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_flavor_s1 AND NOT pio_bitcrusher_flavor_s1_non_bursting_master_requests)))) = '1' then 
        pio_bitcrusher_flavor_s1_slavearbiterlockenable <= or_reduce(pio_bitcrusher_flavor_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_bitcrusher_flavor/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_bitcrusher_flavor_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_bitcrusher_flavor_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_bitcrusher_flavor_s1_slavearbiterlockenable2 <= or_reduce(pio_bitcrusher_flavor_s1_arb_share_counter_next_value);
  --cpu/data_master pio_bitcrusher_flavor/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_bitcrusher_flavor_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_bitcrusher_flavor_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_bitcrusher_flavor_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_flavor_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_bitcrusher_flavor_s1_writedata mux, which is an e_mux
  pio_bitcrusher_flavor_s1_writedata <= cpu_data_master_writedata (3 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_bitcrusher_flavor_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1;
  --cpu/data_master saved-grant pio_bitcrusher_flavor/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_bitcrusher_flavor_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_flavor_s1;
  --allow new arb cycle for pio_bitcrusher_flavor/s1, which is an e_assign
  pio_bitcrusher_flavor_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_bitcrusher_flavor_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_bitcrusher_flavor_s1_master_qreq_vector <= std_logic'('1');
  --pio_bitcrusher_flavor_s1_reset_n assignment, which is an e_assign
  pio_bitcrusher_flavor_s1_reset_n <= reset_n;
  pio_bitcrusher_flavor_s1_chipselect <= internal_cpu_data_master_granted_pio_bitcrusher_flavor_s1;
  --pio_bitcrusher_flavor_s1_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_flavor_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_bitcrusher_flavor_s1_begins_xfer) = '1'), pio_bitcrusher_flavor_s1_unreg_firsttransfer, pio_bitcrusher_flavor_s1_reg_firsttransfer);
  --pio_bitcrusher_flavor_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_flavor_s1_unreg_firsttransfer <= NOT ((pio_bitcrusher_flavor_s1_slavearbiterlockenable AND pio_bitcrusher_flavor_s1_any_continuerequest));
  --pio_bitcrusher_flavor_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_flavor_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_flavor_s1_begins_xfer) = '1' then 
        pio_bitcrusher_flavor_s1_reg_firsttransfer <= pio_bitcrusher_flavor_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_bitcrusher_flavor_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_bitcrusher_flavor_s1_beginbursttransfer_internal <= pio_bitcrusher_flavor_s1_begins_xfer;
  --~pio_bitcrusher_flavor_s1_write_n assignment, which is an e_mux
  pio_bitcrusher_flavor_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_bitcrusher_flavor_s1 AND cpu_data_master_write));
  shifted_address_to_pio_bitcrusher_flavor_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_bitcrusher_flavor_s1_address mux, which is an e_mux
  pio_bitcrusher_flavor_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_bitcrusher_flavor_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_bitcrusher_flavor_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_bitcrusher_flavor_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_bitcrusher_flavor_s1_end_xfer <= pio_bitcrusher_flavor_s1_end_xfer;
    end if;

  end process;

  --pio_bitcrusher_flavor_s1_waits_for_read in a cycle, which is an e_mux
  pio_bitcrusher_flavor_s1_waits_for_read <= pio_bitcrusher_flavor_s1_in_a_read_cycle AND pio_bitcrusher_flavor_s1_begins_xfer;
  --pio_bitcrusher_flavor_s1_in_a_read_cycle assignment, which is an e_assign
  pio_bitcrusher_flavor_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_flavor_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_bitcrusher_flavor_s1_in_a_read_cycle;
  --pio_bitcrusher_flavor_s1_waits_for_write in a cycle, which is an e_mux
  pio_bitcrusher_flavor_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_bitcrusher_flavor_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_bitcrusher_flavor_s1_in_a_write_cycle assignment, which is an e_assign
  pio_bitcrusher_flavor_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_flavor_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_bitcrusher_flavor_s1_in_a_write_cycle;
  wait_for_pio_bitcrusher_flavor_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_bitcrusher_flavor_s1 <= internal_cpu_data_master_granted_pio_bitcrusher_flavor_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_bitcrusher_flavor_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_flavor_s1;
--synthesis translate_off
    --pio_bitcrusher_flavor/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_bitcrusher_tone_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_bitcrusher_tone_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                 signal d1_pio_bitcrusher_tone_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_bitcrusher_tone_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_bitcrusher_tone_s1_chipselect : OUT STD_LOGIC;
                 signal pio_bitcrusher_tone_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_bitcrusher_tone_s1_reset_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_tone_s1_write_n : OUT STD_LOGIC;
                 signal pio_bitcrusher_tone_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_bitcrusher_tone_s1_arbitrator;


architecture europa of pio_bitcrusher_tone_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_allgrants :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_any_continuerequest :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_tone_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_tone_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_bitcrusher_tone_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_begins_xfer :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_end_xfer :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_grant_vector :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_waits_for_read :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_bitcrusher_tone_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_bitcrusher_tone_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_bitcrusher_tone_s1_end_xfer;
    end if;

  end process;

  pio_bitcrusher_tone_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_bitcrusher_tone_s1);
  --assign pio_bitcrusher_tone_s1_readdata_from_sa = pio_bitcrusher_tone_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_bitcrusher_tone_s1_readdata_from_sa <= pio_bitcrusher_tone_s1_readdata;
  internal_cpu_data_master_requests_pio_bitcrusher_tone_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000111000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_bitcrusher_tone_s1_arb_share_counter set values, which is an e_mux
  pio_bitcrusher_tone_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_bitcrusher_tone_s1_non_bursting_master_requests mux, which is an e_mux
  pio_bitcrusher_tone_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_bitcrusher_tone_s1;
  --pio_bitcrusher_tone_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_bitcrusher_tone_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_bitcrusher_tone_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_bitcrusher_tone_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_bitcrusher_tone_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_tone_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_bitcrusher_tone_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_bitcrusher_tone_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_bitcrusher_tone_s1_allgrants all slave grants, which is an e_mux
  pio_bitcrusher_tone_s1_allgrants <= pio_bitcrusher_tone_s1_grant_vector;
  --pio_bitcrusher_tone_s1_end_xfer assignment, which is an e_assign
  pio_bitcrusher_tone_s1_end_xfer <= NOT ((pio_bitcrusher_tone_s1_waits_for_read OR pio_bitcrusher_tone_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_bitcrusher_tone_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_bitcrusher_tone_s1 <= pio_bitcrusher_tone_s1_end_xfer AND (((NOT pio_bitcrusher_tone_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_bitcrusher_tone_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_bitcrusher_tone_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_bitcrusher_tone_s1 AND pio_bitcrusher_tone_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_tone_s1 AND NOT pio_bitcrusher_tone_s1_non_bursting_master_requests));
  --pio_bitcrusher_tone_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_tone_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_tone_s1_arb_counter_enable) = '1' then 
        pio_bitcrusher_tone_s1_arb_share_counter <= pio_bitcrusher_tone_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_bitcrusher_tone_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_tone_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_bitcrusher_tone_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_bitcrusher_tone_s1)) OR ((end_xfer_arb_share_counter_term_pio_bitcrusher_tone_s1 AND NOT pio_bitcrusher_tone_s1_non_bursting_master_requests)))) = '1' then 
        pio_bitcrusher_tone_s1_slavearbiterlockenable <= or_reduce(pio_bitcrusher_tone_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_bitcrusher_tone/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_bitcrusher_tone_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_bitcrusher_tone_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_bitcrusher_tone_s1_slavearbiterlockenable2 <= or_reduce(pio_bitcrusher_tone_s1_arb_share_counter_next_value);
  --cpu/data_master pio_bitcrusher_tone/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_bitcrusher_tone_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_bitcrusher_tone_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_bitcrusher_tone_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_tone_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_bitcrusher_tone_s1_writedata mux, which is an e_mux
  pio_bitcrusher_tone_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_bitcrusher_tone_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_tone_s1;
  --cpu/data_master saved-grant pio_bitcrusher_tone/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_bitcrusher_tone_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_tone_s1;
  --allow new arb cycle for pio_bitcrusher_tone/s1, which is an e_assign
  pio_bitcrusher_tone_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_bitcrusher_tone_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_bitcrusher_tone_s1_master_qreq_vector <= std_logic'('1');
  --pio_bitcrusher_tone_s1_reset_n assignment, which is an e_assign
  pio_bitcrusher_tone_s1_reset_n <= reset_n;
  pio_bitcrusher_tone_s1_chipselect <= internal_cpu_data_master_granted_pio_bitcrusher_tone_s1;
  --pio_bitcrusher_tone_s1_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_tone_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_bitcrusher_tone_s1_begins_xfer) = '1'), pio_bitcrusher_tone_s1_unreg_firsttransfer, pio_bitcrusher_tone_s1_reg_firsttransfer);
  --pio_bitcrusher_tone_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_bitcrusher_tone_s1_unreg_firsttransfer <= NOT ((pio_bitcrusher_tone_s1_slavearbiterlockenable AND pio_bitcrusher_tone_s1_any_continuerequest));
  --pio_bitcrusher_tone_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_bitcrusher_tone_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_bitcrusher_tone_s1_begins_xfer) = '1' then 
        pio_bitcrusher_tone_s1_reg_firsttransfer <= pio_bitcrusher_tone_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_bitcrusher_tone_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_bitcrusher_tone_s1_beginbursttransfer_internal <= pio_bitcrusher_tone_s1_begins_xfer;
  --~pio_bitcrusher_tone_s1_write_n assignment, which is an e_mux
  pio_bitcrusher_tone_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_bitcrusher_tone_s1 AND cpu_data_master_write));
  shifted_address_to_pio_bitcrusher_tone_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_bitcrusher_tone_s1_address mux, which is an e_mux
  pio_bitcrusher_tone_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_bitcrusher_tone_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_bitcrusher_tone_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_bitcrusher_tone_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_bitcrusher_tone_s1_end_xfer <= pio_bitcrusher_tone_s1_end_xfer;
    end if;

  end process;

  --pio_bitcrusher_tone_s1_waits_for_read in a cycle, which is an e_mux
  pio_bitcrusher_tone_s1_waits_for_read <= pio_bitcrusher_tone_s1_in_a_read_cycle AND pio_bitcrusher_tone_s1_begins_xfer;
  --pio_bitcrusher_tone_s1_in_a_read_cycle assignment, which is an e_assign
  pio_bitcrusher_tone_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_tone_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_bitcrusher_tone_s1_in_a_read_cycle;
  --pio_bitcrusher_tone_s1_waits_for_write in a cycle, which is an e_mux
  pio_bitcrusher_tone_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_bitcrusher_tone_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_bitcrusher_tone_s1_in_a_write_cycle assignment, which is an e_assign
  pio_bitcrusher_tone_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_bitcrusher_tone_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_bitcrusher_tone_s1_in_a_write_cycle;
  wait_for_pio_bitcrusher_tone_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_bitcrusher_tone_s1 <= internal_cpu_data_master_granted_pio_bitcrusher_tone_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 <= internal_cpu_data_master_qualified_request_pio_bitcrusher_tone_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_bitcrusher_tone_s1 <= internal_cpu_data_master_requests_pio_bitcrusher_tone_s1;
--synthesis translate_off
    --pio_bitcrusher_tone/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_compressor_bypass_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_compressor_bypass_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                 signal d1_pio_compressor_bypass_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_compressor_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_compressor_bypass_s1_chipselect : OUT STD_LOGIC;
                 signal pio_compressor_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_compressor_bypass_s1_reset_n : OUT STD_LOGIC;
                 signal pio_compressor_bypass_s1_write_n : OUT STD_LOGIC;
                 signal pio_compressor_bypass_s1_writedata : OUT STD_LOGIC
              );
end entity pio_compressor_bypass_s1_arbitrator;


architecture europa of pio_compressor_bypass_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal pio_compressor_bypass_s1_allgrants :  STD_LOGIC;
                signal pio_compressor_bypass_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_compressor_bypass_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_compressor_bypass_s1_any_continuerequest :  STD_LOGIC;
                signal pio_compressor_bypass_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_compressor_bypass_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_bypass_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_bypass_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_bypass_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_compressor_bypass_s1_begins_xfer :  STD_LOGIC;
                signal pio_compressor_bypass_s1_end_xfer :  STD_LOGIC;
                signal pio_compressor_bypass_s1_firsttransfer :  STD_LOGIC;
                signal pio_compressor_bypass_s1_grant_vector :  STD_LOGIC;
                signal pio_compressor_bypass_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_compressor_bypass_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_compressor_bypass_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_compressor_bypass_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_compressor_bypass_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_compressor_bypass_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_compressor_bypass_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_compressor_bypass_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_compressor_bypass_s1_waits_for_read :  STD_LOGIC;
                signal pio_compressor_bypass_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_compressor_bypass_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_compressor_bypass_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_compressor_bypass_s1_end_xfer;
    end if;

  end process;

  pio_compressor_bypass_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_compressor_bypass_s1);
  --assign pio_compressor_bypass_s1_readdata_from_sa = pio_compressor_bypass_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_compressor_bypass_s1_readdata_from_sa <= pio_compressor_bypass_s1_readdata;
  internal_cpu_data_master_requests_pio_compressor_bypass_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000011100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_compressor_bypass_s1_arb_share_counter set values, which is an e_mux
  pio_compressor_bypass_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_compressor_bypass_s1_non_bursting_master_requests mux, which is an e_mux
  pio_compressor_bypass_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_compressor_bypass_s1;
  --pio_compressor_bypass_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_compressor_bypass_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_compressor_bypass_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_compressor_bypass_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_compressor_bypass_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_compressor_bypass_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_compressor_bypass_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_compressor_bypass_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_compressor_bypass_s1_allgrants all slave grants, which is an e_mux
  pio_compressor_bypass_s1_allgrants <= pio_compressor_bypass_s1_grant_vector;
  --pio_compressor_bypass_s1_end_xfer assignment, which is an e_assign
  pio_compressor_bypass_s1_end_xfer <= NOT ((pio_compressor_bypass_s1_waits_for_read OR pio_compressor_bypass_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_compressor_bypass_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_compressor_bypass_s1 <= pio_compressor_bypass_s1_end_xfer AND (((NOT pio_compressor_bypass_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_compressor_bypass_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_compressor_bypass_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_compressor_bypass_s1 AND pio_compressor_bypass_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_compressor_bypass_s1 AND NOT pio_compressor_bypass_s1_non_bursting_master_requests));
  --pio_compressor_bypass_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_bypass_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_compressor_bypass_s1_arb_counter_enable) = '1' then 
        pio_compressor_bypass_s1_arb_share_counter <= pio_compressor_bypass_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_compressor_bypass_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_bypass_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_compressor_bypass_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_compressor_bypass_s1)) OR ((end_xfer_arb_share_counter_term_pio_compressor_bypass_s1 AND NOT pio_compressor_bypass_s1_non_bursting_master_requests)))) = '1' then 
        pio_compressor_bypass_s1_slavearbiterlockenable <= or_reduce(pio_compressor_bypass_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_compressor_bypass/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_compressor_bypass_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_compressor_bypass_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_compressor_bypass_s1_slavearbiterlockenable2 <= or_reduce(pio_compressor_bypass_s1_arb_share_counter_next_value);
  --cpu/data_master pio_compressor_bypass/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_compressor_bypass_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_compressor_bypass_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_compressor_bypass_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_compressor_bypass_s1 <= internal_cpu_data_master_requests_pio_compressor_bypass_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_compressor_bypass_s1_writedata mux, which is an e_mux
  pio_compressor_bypass_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_compressor_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_compressor_bypass_s1;
  --cpu/data_master saved-grant pio_compressor_bypass/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_compressor_bypass_s1 <= internal_cpu_data_master_requests_pio_compressor_bypass_s1;
  --allow new arb cycle for pio_compressor_bypass/s1, which is an e_assign
  pio_compressor_bypass_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_compressor_bypass_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_compressor_bypass_s1_master_qreq_vector <= std_logic'('1');
  --pio_compressor_bypass_s1_reset_n assignment, which is an e_assign
  pio_compressor_bypass_s1_reset_n <= reset_n;
  pio_compressor_bypass_s1_chipselect <= internal_cpu_data_master_granted_pio_compressor_bypass_s1;
  --pio_compressor_bypass_s1_firsttransfer first transaction, which is an e_assign
  pio_compressor_bypass_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_compressor_bypass_s1_begins_xfer) = '1'), pio_compressor_bypass_s1_unreg_firsttransfer, pio_compressor_bypass_s1_reg_firsttransfer);
  --pio_compressor_bypass_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_compressor_bypass_s1_unreg_firsttransfer <= NOT ((pio_compressor_bypass_s1_slavearbiterlockenable AND pio_compressor_bypass_s1_any_continuerequest));
  --pio_compressor_bypass_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_bypass_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_compressor_bypass_s1_begins_xfer) = '1' then 
        pio_compressor_bypass_s1_reg_firsttransfer <= pio_compressor_bypass_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_compressor_bypass_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_compressor_bypass_s1_beginbursttransfer_internal <= pio_compressor_bypass_s1_begins_xfer;
  --~pio_compressor_bypass_s1_write_n assignment, which is an e_mux
  pio_compressor_bypass_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_compressor_bypass_s1 AND cpu_data_master_write));
  shifted_address_to_pio_compressor_bypass_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_compressor_bypass_s1_address mux, which is an e_mux
  pio_compressor_bypass_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_compressor_bypass_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_compressor_bypass_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_compressor_bypass_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_compressor_bypass_s1_end_xfer <= pio_compressor_bypass_s1_end_xfer;
    end if;

  end process;

  --pio_compressor_bypass_s1_waits_for_read in a cycle, which is an e_mux
  pio_compressor_bypass_s1_waits_for_read <= pio_compressor_bypass_s1_in_a_read_cycle AND pio_compressor_bypass_s1_begins_xfer;
  --pio_compressor_bypass_s1_in_a_read_cycle assignment, which is an e_assign
  pio_compressor_bypass_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_compressor_bypass_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_compressor_bypass_s1_in_a_read_cycle;
  --pio_compressor_bypass_s1_waits_for_write in a cycle, which is an e_mux
  pio_compressor_bypass_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_compressor_bypass_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_compressor_bypass_s1_in_a_write_cycle assignment, which is an e_assign
  pio_compressor_bypass_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_compressor_bypass_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_compressor_bypass_s1_in_a_write_cycle;
  wait_for_pio_compressor_bypass_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_compressor_bypass_s1 <= internal_cpu_data_master_granted_pio_compressor_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_compressor_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_compressor_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_compressor_bypass_s1 <= internal_cpu_data_master_requests_pio_compressor_bypass_s1;
--synthesis translate_off
    --pio_compressor_bypass/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_compressor_gain_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_compressor_gain_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_compressor_gain_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_compressor_gain_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_compressor_gain_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_compressor_gain_s1 : OUT STD_LOGIC;
                 signal d1_pio_compressor_gain_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_compressor_gain_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_compressor_gain_s1_chipselect : OUT STD_LOGIC;
                 signal pio_compressor_gain_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pio_compressor_gain_s1_reset_n : OUT STD_LOGIC;
                 signal pio_compressor_gain_s1_write_n : OUT STD_LOGIC;
                 signal pio_compressor_gain_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity pio_compressor_gain_s1_arbitrator;


architecture europa of pio_compressor_gain_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_compressor_gain_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_compressor_gain_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_compressor_gain_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_compressor_gain_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_compressor_gain_s1 :  STD_LOGIC;
                signal pio_compressor_gain_s1_allgrants :  STD_LOGIC;
                signal pio_compressor_gain_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_compressor_gain_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_compressor_gain_s1_any_continuerequest :  STD_LOGIC;
                signal pio_compressor_gain_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_compressor_gain_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_gain_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_gain_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_gain_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_compressor_gain_s1_begins_xfer :  STD_LOGIC;
                signal pio_compressor_gain_s1_end_xfer :  STD_LOGIC;
                signal pio_compressor_gain_s1_firsttransfer :  STD_LOGIC;
                signal pio_compressor_gain_s1_grant_vector :  STD_LOGIC;
                signal pio_compressor_gain_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_compressor_gain_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_compressor_gain_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_compressor_gain_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_compressor_gain_s1_pretend_byte_enable :  STD_LOGIC;
                signal pio_compressor_gain_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_compressor_gain_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_compressor_gain_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_compressor_gain_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_compressor_gain_s1_waits_for_read :  STD_LOGIC;
                signal pio_compressor_gain_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_compressor_gain_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_compressor_gain_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_compressor_gain_s1_end_xfer;
    end if;

  end process;

  pio_compressor_gain_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_compressor_gain_s1);
  --assign pio_compressor_gain_s1_readdata_from_sa = pio_compressor_gain_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_compressor_gain_s1_readdata_from_sa <= pio_compressor_gain_s1_readdata;
  internal_cpu_data_master_requests_pio_compressor_gain_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000011000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_compressor_gain_s1_arb_share_counter set values, which is an e_mux
  pio_compressor_gain_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_compressor_gain_s1_non_bursting_master_requests mux, which is an e_mux
  pio_compressor_gain_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_compressor_gain_s1;
  --pio_compressor_gain_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_compressor_gain_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_compressor_gain_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_compressor_gain_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_compressor_gain_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_compressor_gain_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_compressor_gain_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_compressor_gain_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_compressor_gain_s1_allgrants all slave grants, which is an e_mux
  pio_compressor_gain_s1_allgrants <= pio_compressor_gain_s1_grant_vector;
  --pio_compressor_gain_s1_end_xfer assignment, which is an e_assign
  pio_compressor_gain_s1_end_xfer <= NOT ((pio_compressor_gain_s1_waits_for_read OR pio_compressor_gain_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_compressor_gain_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_compressor_gain_s1 <= pio_compressor_gain_s1_end_xfer AND (((NOT pio_compressor_gain_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_compressor_gain_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_compressor_gain_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_compressor_gain_s1 AND pio_compressor_gain_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_compressor_gain_s1 AND NOT pio_compressor_gain_s1_non_bursting_master_requests));
  --pio_compressor_gain_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_gain_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_compressor_gain_s1_arb_counter_enable) = '1' then 
        pio_compressor_gain_s1_arb_share_counter <= pio_compressor_gain_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_compressor_gain_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_gain_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_compressor_gain_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_compressor_gain_s1)) OR ((end_xfer_arb_share_counter_term_pio_compressor_gain_s1 AND NOT pio_compressor_gain_s1_non_bursting_master_requests)))) = '1' then 
        pio_compressor_gain_s1_slavearbiterlockenable <= or_reduce(pio_compressor_gain_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_compressor_gain/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_compressor_gain_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_compressor_gain_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_compressor_gain_s1_slavearbiterlockenable2 <= or_reduce(pio_compressor_gain_s1_arb_share_counter_next_value);
  --cpu/data_master pio_compressor_gain/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_compressor_gain_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_compressor_gain_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_compressor_gain_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_compressor_gain_s1 <= internal_cpu_data_master_requests_pio_compressor_gain_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_compressor_gain_s1_writedata mux, which is an e_mux
  pio_compressor_gain_s1_writedata <= cpu_data_master_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_compressor_gain_s1 <= internal_cpu_data_master_qualified_request_pio_compressor_gain_s1;
  --cpu/data_master saved-grant pio_compressor_gain/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_compressor_gain_s1 <= internal_cpu_data_master_requests_pio_compressor_gain_s1;
  --allow new arb cycle for pio_compressor_gain/s1, which is an e_assign
  pio_compressor_gain_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_compressor_gain_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_compressor_gain_s1_master_qreq_vector <= std_logic'('1');
  --pio_compressor_gain_s1_reset_n assignment, which is an e_assign
  pio_compressor_gain_s1_reset_n <= reset_n;
  pio_compressor_gain_s1_chipselect <= internal_cpu_data_master_granted_pio_compressor_gain_s1;
  --pio_compressor_gain_s1_firsttransfer first transaction, which is an e_assign
  pio_compressor_gain_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_compressor_gain_s1_begins_xfer) = '1'), pio_compressor_gain_s1_unreg_firsttransfer, pio_compressor_gain_s1_reg_firsttransfer);
  --pio_compressor_gain_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_compressor_gain_s1_unreg_firsttransfer <= NOT ((pio_compressor_gain_s1_slavearbiterlockenable AND pio_compressor_gain_s1_any_continuerequest));
  --pio_compressor_gain_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_gain_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_compressor_gain_s1_begins_xfer) = '1' then 
        pio_compressor_gain_s1_reg_firsttransfer <= pio_compressor_gain_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_compressor_gain_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_compressor_gain_s1_beginbursttransfer_internal <= pio_compressor_gain_s1_begins_xfer;
  --~pio_compressor_gain_s1_write_n assignment, which is an e_mux
  pio_compressor_gain_s1_write_n <= NOT ((((internal_cpu_data_master_granted_pio_compressor_gain_s1 AND cpu_data_master_write)) AND pio_compressor_gain_s1_pretend_byte_enable));
  shifted_address_to_pio_compressor_gain_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_compressor_gain_s1_address mux, which is an e_mux
  pio_compressor_gain_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_compressor_gain_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_compressor_gain_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_compressor_gain_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_compressor_gain_s1_end_xfer <= pio_compressor_gain_s1_end_xfer;
    end if;

  end process;

  --pio_compressor_gain_s1_waits_for_read in a cycle, which is an e_mux
  pio_compressor_gain_s1_waits_for_read <= pio_compressor_gain_s1_in_a_read_cycle AND pio_compressor_gain_s1_begins_xfer;
  --pio_compressor_gain_s1_in_a_read_cycle assignment, which is an e_assign
  pio_compressor_gain_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_compressor_gain_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_compressor_gain_s1_in_a_read_cycle;
  --pio_compressor_gain_s1_waits_for_write in a cycle, which is an e_mux
  pio_compressor_gain_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_compressor_gain_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_compressor_gain_s1_in_a_write_cycle assignment, which is an e_assign
  pio_compressor_gain_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_compressor_gain_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_compressor_gain_s1_in_a_write_cycle;
  wait_for_pio_compressor_gain_s1_counter <= std_logic'('0');
  --pio_compressor_gain_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  pio_compressor_gain_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pio_compressor_gain_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_compressor_gain_s1 <= internal_cpu_data_master_granted_pio_compressor_gain_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_compressor_gain_s1 <= internal_cpu_data_master_qualified_request_pio_compressor_gain_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_compressor_gain_s1 <= internal_cpu_data_master_requests_pio_compressor_gain_s1;
--synthesis translate_off
    --pio_compressor_gain/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_compressor_treshold_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_compressor_treshold_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                 signal d1_pio_compressor_treshold_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_compressor_treshold_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_compressor_treshold_s1_chipselect : OUT STD_LOGIC;
                 signal pio_compressor_treshold_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_compressor_treshold_s1_reset_n : OUT STD_LOGIC;
                 signal pio_compressor_treshold_s1_write_n : OUT STD_LOGIC;
                 signal pio_compressor_treshold_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_compressor_treshold_s1_arbitrator;


architecture europa of pio_compressor_treshold_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal pio_compressor_treshold_s1_allgrants :  STD_LOGIC;
                signal pio_compressor_treshold_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_compressor_treshold_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_compressor_treshold_s1_any_continuerequest :  STD_LOGIC;
                signal pio_compressor_treshold_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_compressor_treshold_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_treshold_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_treshold_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_compressor_treshold_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_compressor_treshold_s1_begins_xfer :  STD_LOGIC;
                signal pio_compressor_treshold_s1_end_xfer :  STD_LOGIC;
                signal pio_compressor_treshold_s1_firsttransfer :  STD_LOGIC;
                signal pio_compressor_treshold_s1_grant_vector :  STD_LOGIC;
                signal pio_compressor_treshold_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_compressor_treshold_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_compressor_treshold_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_compressor_treshold_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_compressor_treshold_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_compressor_treshold_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_compressor_treshold_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_compressor_treshold_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_compressor_treshold_s1_waits_for_read :  STD_LOGIC;
                signal pio_compressor_treshold_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_compressor_treshold_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_compressor_treshold_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_compressor_treshold_s1_end_xfer;
    end if;

  end process;

  pio_compressor_treshold_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_compressor_treshold_s1);
  --assign pio_compressor_treshold_s1_readdata_from_sa = pio_compressor_treshold_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_compressor_treshold_s1_readdata_from_sa <= pio_compressor_treshold_s1_readdata;
  internal_cpu_data_master_requests_pio_compressor_treshold_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000011010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_compressor_treshold_s1_arb_share_counter set values, which is an e_mux
  pio_compressor_treshold_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_compressor_treshold_s1_non_bursting_master_requests mux, which is an e_mux
  pio_compressor_treshold_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_compressor_treshold_s1;
  --pio_compressor_treshold_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_compressor_treshold_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_compressor_treshold_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_compressor_treshold_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_compressor_treshold_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_compressor_treshold_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_compressor_treshold_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_compressor_treshold_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_compressor_treshold_s1_allgrants all slave grants, which is an e_mux
  pio_compressor_treshold_s1_allgrants <= pio_compressor_treshold_s1_grant_vector;
  --pio_compressor_treshold_s1_end_xfer assignment, which is an e_assign
  pio_compressor_treshold_s1_end_xfer <= NOT ((pio_compressor_treshold_s1_waits_for_read OR pio_compressor_treshold_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_compressor_treshold_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_compressor_treshold_s1 <= pio_compressor_treshold_s1_end_xfer AND (((NOT pio_compressor_treshold_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_compressor_treshold_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_compressor_treshold_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_compressor_treshold_s1 AND pio_compressor_treshold_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_compressor_treshold_s1 AND NOT pio_compressor_treshold_s1_non_bursting_master_requests));
  --pio_compressor_treshold_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_treshold_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_compressor_treshold_s1_arb_counter_enable) = '1' then 
        pio_compressor_treshold_s1_arb_share_counter <= pio_compressor_treshold_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_compressor_treshold_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_treshold_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_compressor_treshold_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_compressor_treshold_s1)) OR ((end_xfer_arb_share_counter_term_pio_compressor_treshold_s1 AND NOT pio_compressor_treshold_s1_non_bursting_master_requests)))) = '1' then 
        pio_compressor_treshold_s1_slavearbiterlockenable <= or_reduce(pio_compressor_treshold_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_compressor_treshold/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_compressor_treshold_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_compressor_treshold_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_compressor_treshold_s1_slavearbiterlockenable2 <= or_reduce(pio_compressor_treshold_s1_arb_share_counter_next_value);
  --cpu/data_master pio_compressor_treshold/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_compressor_treshold_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_compressor_treshold_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_compressor_treshold_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_compressor_treshold_s1 <= internal_cpu_data_master_requests_pio_compressor_treshold_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_compressor_treshold_s1_writedata mux, which is an e_mux
  pio_compressor_treshold_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_compressor_treshold_s1 <= internal_cpu_data_master_qualified_request_pio_compressor_treshold_s1;
  --cpu/data_master saved-grant pio_compressor_treshold/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_compressor_treshold_s1 <= internal_cpu_data_master_requests_pio_compressor_treshold_s1;
  --allow new arb cycle for pio_compressor_treshold/s1, which is an e_assign
  pio_compressor_treshold_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_compressor_treshold_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_compressor_treshold_s1_master_qreq_vector <= std_logic'('1');
  --pio_compressor_treshold_s1_reset_n assignment, which is an e_assign
  pio_compressor_treshold_s1_reset_n <= reset_n;
  pio_compressor_treshold_s1_chipselect <= internal_cpu_data_master_granted_pio_compressor_treshold_s1;
  --pio_compressor_treshold_s1_firsttransfer first transaction, which is an e_assign
  pio_compressor_treshold_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_compressor_treshold_s1_begins_xfer) = '1'), pio_compressor_treshold_s1_unreg_firsttransfer, pio_compressor_treshold_s1_reg_firsttransfer);
  --pio_compressor_treshold_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_compressor_treshold_s1_unreg_firsttransfer <= NOT ((pio_compressor_treshold_s1_slavearbiterlockenable AND pio_compressor_treshold_s1_any_continuerequest));
  --pio_compressor_treshold_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_compressor_treshold_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_compressor_treshold_s1_begins_xfer) = '1' then 
        pio_compressor_treshold_s1_reg_firsttransfer <= pio_compressor_treshold_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_compressor_treshold_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_compressor_treshold_s1_beginbursttransfer_internal <= pio_compressor_treshold_s1_begins_xfer;
  --~pio_compressor_treshold_s1_write_n assignment, which is an e_mux
  pio_compressor_treshold_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_compressor_treshold_s1 AND cpu_data_master_write));
  shifted_address_to_pio_compressor_treshold_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_compressor_treshold_s1_address mux, which is an e_mux
  pio_compressor_treshold_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_compressor_treshold_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_compressor_treshold_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_compressor_treshold_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_compressor_treshold_s1_end_xfer <= pio_compressor_treshold_s1_end_xfer;
    end if;

  end process;

  --pio_compressor_treshold_s1_waits_for_read in a cycle, which is an e_mux
  pio_compressor_treshold_s1_waits_for_read <= pio_compressor_treshold_s1_in_a_read_cycle AND pio_compressor_treshold_s1_begins_xfer;
  --pio_compressor_treshold_s1_in_a_read_cycle assignment, which is an e_assign
  pio_compressor_treshold_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_compressor_treshold_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_compressor_treshold_s1_in_a_read_cycle;
  --pio_compressor_treshold_s1_waits_for_write in a cycle, which is an e_mux
  pio_compressor_treshold_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_compressor_treshold_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_compressor_treshold_s1_in_a_write_cycle assignment, which is an e_assign
  pio_compressor_treshold_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_compressor_treshold_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_compressor_treshold_s1_in_a_write_cycle;
  wait_for_pio_compressor_treshold_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_compressor_treshold_s1 <= internal_cpu_data_master_granted_pio_compressor_treshold_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_compressor_treshold_s1 <= internal_cpu_data_master_qualified_request_pio_compressor_treshold_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_compressor_treshold_s1 <= internal_cpu_data_master_requests_pio_compressor_treshold_s1;
--synthesis translate_off
    --pio_compressor_treshold/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_delay_bypass_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_delay_bypass_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_delay_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_delay_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_delay_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_delay_bypass_s1 : OUT STD_LOGIC;
                 signal d1_pio_delay_bypass_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_delay_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_delay_bypass_s1_chipselect : OUT STD_LOGIC;
                 signal pio_delay_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_delay_bypass_s1_reset_n : OUT STD_LOGIC;
                 signal pio_delay_bypass_s1_write_n : OUT STD_LOGIC;
                 signal pio_delay_bypass_s1_writedata : OUT STD_LOGIC
              );
end entity pio_delay_bypass_s1_arbitrator;


architecture europa of pio_delay_bypass_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_delay_bypass_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_delay_bypass_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_delay_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_delay_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_delay_bypass_s1 :  STD_LOGIC;
                signal pio_delay_bypass_s1_allgrants :  STD_LOGIC;
                signal pio_delay_bypass_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_delay_bypass_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_delay_bypass_s1_any_continuerequest :  STD_LOGIC;
                signal pio_delay_bypass_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_delay_bypass_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_bypass_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_bypass_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_bypass_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_delay_bypass_s1_begins_xfer :  STD_LOGIC;
                signal pio_delay_bypass_s1_end_xfer :  STD_LOGIC;
                signal pio_delay_bypass_s1_firsttransfer :  STD_LOGIC;
                signal pio_delay_bypass_s1_grant_vector :  STD_LOGIC;
                signal pio_delay_bypass_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_delay_bypass_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_delay_bypass_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_delay_bypass_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_delay_bypass_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_delay_bypass_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_delay_bypass_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_delay_bypass_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_delay_bypass_s1_waits_for_read :  STD_LOGIC;
                signal pio_delay_bypass_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_delay_bypass_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_delay_bypass_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_delay_bypass_s1_end_xfer;
    end if;

  end process;

  pio_delay_bypass_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_delay_bypass_s1);
  --assign pio_delay_bypass_s1_readdata_from_sa = pio_delay_bypass_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_delay_bypass_s1_readdata_from_sa <= pio_delay_bypass_s1_readdata;
  internal_cpu_data_master_requests_pio_delay_bypass_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000001010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_delay_bypass_s1_arb_share_counter set values, which is an e_mux
  pio_delay_bypass_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_delay_bypass_s1_non_bursting_master_requests mux, which is an e_mux
  pio_delay_bypass_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_delay_bypass_s1;
  --pio_delay_bypass_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_delay_bypass_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_delay_bypass_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_delay_bypass_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_delay_bypass_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_delay_bypass_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_delay_bypass_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_delay_bypass_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_delay_bypass_s1_allgrants all slave grants, which is an e_mux
  pio_delay_bypass_s1_allgrants <= pio_delay_bypass_s1_grant_vector;
  --pio_delay_bypass_s1_end_xfer assignment, which is an e_assign
  pio_delay_bypass_s1_end_xfer <= NOT ((pio_delay_bypass_s1_waits_for_read OR pio_delay_bypass_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_delay_bypass_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_delay_bypass_s1 <= pio_delay_bypass_s1_end_xfer AND (((NOT pio_delay_bypass_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_delay_bypass_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_delay_bypass_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_delay_bypass_s1 AND pio_delay_bypass_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_delay_bypass_s1 AND NOT pio_delay_bypass_s1_non_bursting_master_requests));
  --pio_delay_bypass_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_bypass_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_delay_bypass_s1_arb_counter_enable) = '1' then 
        pio_delay_bypass_s1_arb_share_counter <= pio_delay_bypass_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_delay_bypass_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_bypass_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_delay_bypass_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_delay_bypass_s1)) OR ((end_xfer_arb_share_counter_term_pio_delay_bypass_s1 AND NOT pio_delay_bypass_s1_non_bursting_master_requests)))) = '1' then 
        pio_delay_bypass_s1_slavearbiterlockenable <= or_reduce(pio_delay_bypass_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_delay_bypass/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_delay_bypass_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_delay_bypass_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_delay_bypass_s1_slavearbiterlockenable2 <= or_reduce(pio_delay_bypass_s1_arb_share_counter_next_value);
  --cpu/data_master pio_delay_bypass/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_delay_bypass_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_delay_bypass_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_delay_bypass_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_delay_bypass_s1 <= internal_cpu_data_master_requests_pio_delay_bypass_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_delay_bypass_s1_writedata mux, which is an e_mux
  pio_delay_bypass_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_delay_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_delay_bypass_s1;
  --cpu/data_master saved-grant pio_delay_bypass/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_delay_bypass_s1 <= internal_cpu_data_master_requests_pio_delay_bypass_s1;
  --allow new arb cycle for pio_delay_bypass/s1, which is an e_assign
  pio_delay_bypass_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_delay_bypass_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_delay_bypass_s1_master_qreq_vector <= std_logic'('1');
  --pio_delay_bypass_s1_reset_n assignment, which is an e_assign
  pio_delay_bypass_s1_reset_n <= reset_n;
  pio_delay_bypass_s1_chipselect <= internal_cpu_data_master_granted_pio_delay_bypass_s1;
  --pio_delay_bypass_s1_firsttransfer first transaction, which is an e_assign
  pio_delay_bypass_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_delay_bypass_s1_begins_xfer) = '1'), pio_delay_bypass_s1_unreg_firsttransfer, pio_delay_bypass_s1_reg_firsttransfer);
  --pio_delay_bypass_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_delay_bypass_s1_unreg_firsttransfer <= NOT ((pio_delay_bypass_s1_slavearbiterlockenable AND pio_delay_bypass_s1_any_continuerequest));
  --pio_delay_bypass_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_bypass_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_delay_bypass_s1_begins_xfer) = '1' then 
        pio_delay_bypass_s1_reg_firsttransfer <= pio_delay_bypass_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_delay_bypass_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_delay_bypass_s1_beginbursttransfer_internal <= pio_delay_bypass_s1_begins_xfer;
  --~pio_delay_bypass_s1_write_n assignment, which is an e_mux
  pio_delay_bypass_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_delay_bypass_s1 AND cpu_data_master_write));
  shifted_address_to_pio_delay_bypass_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_delay_bypass_s1_address mux, which is an e_mux
  pio_delay_bypass_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_delay_bypass_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_delay_bypass_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_delay_bypass_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_delay_bypass_s1_end_xfer <= pio_delay_bypass_s1_end_xfer;
    end if;

  end process;

  --pio_delay_bypass_s1_waits_for_read in a cycle, which is an e_mux
  pio_delay_bypass_s1_waits_for_read <= pio_delay_bypass_s1_in_a_read_cycle AND pio_delay_bypass_s1_begins_xfer;
  --pio_delay_bypass_s1_in_a_read_cycle assignment, which is an e_assign
  pio_delay_bypass_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_delay_bypass_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_delay_bypass_s1_in_a_read_cycle;
  --pio_delay_bypass_s1_waits_for_write in a cycle, which is an e_mux
  pio_delay_bypass_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_delay_bypass_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_delay_bypass_s1_in_a_write_cycle assignment, which is an e_assign
  pio_delay_bypass_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_delay_bypass_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_delay_bypass_s1_in_a_write_cycle;
  wait_for_pio_delay_bypass_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_delay_bypass_s1 <= internal_cpu_data_master_granted_pio_delay_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_delay_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_delay_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_delay_bypass_s1 <= internal_cpu_data_master_requests_pio_delay_bypass_s1;
--synthesis translate_off
    --pio_delay_bypass/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_delay_decay_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_delay_decay_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_delay_decay_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_delay_decay_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_delay_decay_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_delay_decay_s1 : OUT STD_LOGIC;
                 signal d1_pio_delay_decay_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_delay_decay_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_delay_decay_s1_chipselect : OUT STD_LOGIC;
                 signal pio_delay_decay_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pio_delay_decay_s1_reset_n : OUT STD_LOGIC;
                 signal pio_delay_decay_s1_write_n : OUT STD_LOGIC;
                 signal pio_delay_decay_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity pio_delay_decay_s1_arbitrator;


architecture europa of pio_delay_decay_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_delay_decay_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_delay_decay_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_delay_decay_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_delay_decay_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_delay_decay_s1 :  STD_LOGIC;
                signal pio_delay_decay_s1_allgrants :  STD_LOGIC;
                signal pio_delay_decay_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_delay_decay_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_delay_decay_s1_any_continuerequest :  STD_LOGIC;
                signal pio_delay_decay_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_delay_decay_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_decay_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_decay_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_decay_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_delay_decay_s1_begins_xfer :  STD_LOGIC;
                signal pio_delay_decay_s1_end_xfer :  STD_LOGIC;
                signal pio_delay_decay_s1_firsttransfer :  STD_LOGIC;
                signal pio_delay_decay_s1_grant_vector :  STD_LOGIC;
                signal pio_delay_decay_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_delay_decay_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_delay_decay_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_delay_decay_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_delay_decay_s1_pretend_byte_enable :  STD_LOGIC;
                signal pio_delay_decay_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_delay_decay_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_delay_decay_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_delay_decay_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_delay_decay_s1_waits_for_read :  STD_LOGIC;
                signal pio_delay_decay_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_delay_decay_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_delay_decay_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_delay_decay_s1_end_xfer;
    end if;

  end process;

  pio_delay_decay_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_delay_decay_s1);
  --assign pio_delay_decay_s1_readdata_from_sa = pio_delay_decay_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_delay_decay_s1_readdata_from_sa <= pio_delay_decay_s1_readdata;
  internal_cpu_data_master_requests_pio_delay_decay_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000010000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_delay_decay_s1_arb_share_counter set values, which is an e_mux
  pio_delay_decay_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_delay_decay_s1_non_bursting_master_requests mux, which is an e_mux
  pio_delay_decay_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_delay_decay_s1;
  --pio_delay_decay_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_delay_decay_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_delay_decay_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_delay_decay_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_delay_decay_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_delay_decay_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_delay_decay_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_delay_decay_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_delay_decay_s1_allgrants all slave grants, which is an e_mux
  pio_delay_decay_s1_allgrants <= pio_delay_decay_s1_grant_vector;
  --pio_delay_decay_s1_end_xfer assignment, which is an e_assign
  pio_delay_decay_s1_end_xfer <= NOT ((pio_delay_decay_s1_waits_for_read OR pio_delay_decay_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_delay_decay_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_delay_decay_s1 <= pio_delay_decay_s1_end_xfer AND (((NOT pio_delay_decay_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_delay_decay_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_delay_decay_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_delay_decay_s1 AND pio_delay_decay_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_delay_decay_s1 AND NOT pio_delay_decay_s1_non_bursting_master_requests));
  --pio_delay_decay_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_decay_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_delay_decay_s1_arb_counter_enable) = '1' then 
        pio_delay_decay_s1_arb_share_counter <= pio_delay_decay_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_delay_decay_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_decay_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_delay_decay_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_delay_decay_s1)) OR ((end_xfer_arb_share_counter_term_pio_delay_decay_s1 AND NOT pio_delay_decay_s1_non_bursting_master_requests)))) = '1' then 
        pio_delay_decay_s1_slavearbiterlockenable <= or_reduce(pio_delay_decay_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_delay_decay/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_delay_decay_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_delay_decay_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_delay_decay_s1_slavearbiterlockenable2 <= or_reduce(pio_delay_decay_s1_arb_share_counter_next_value);
  --cpu/data_master pio_delay_decay/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_delay_decay_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_delay_decay_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_delay_decay_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_delay_decay_s1 <= internal_cpu_data_master_requests_pio_delay_decay_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_delay_decay_s1_writedata mux, which is an e_mux
  pio_delay_decay_s1_writedata <= cpu_data_master_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_delay_decay_s1 <= internal_cpu_data_master_qualified_request_pio_delay_decay_s1;
  --cpu/data_master saved-grant pio_delay_decay/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_delay_decay_s1 <= internal_cpu_data_master_requests_pio_delay_decay_s1;
  --allow new arb cycle for pio_delay_decay/s1, which is an e_assign
  pio_delay_decay_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_delay_decay_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_delay_decay_s1_master_qreq_vector <= std_logic'('1');
  --pio_delay_decay_s1_reset_n assignment, which is an e_assign
  pio_delay_decay_s1_reset_n <= reset_n;
  pio_delay_decay_s1_chipselect <= internal_cpu_data_master_granted_pio_delay_decay_s1;
  --pio_delay_decay_s1_firsttransfer first transaction, which is an e_assign
  pio_delay_decay_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_delay_decay_s1_begins_xfer) = '1'), pio_delay_decay_s1_unreg_firsttransfer, pio_delay_decay_s1_reg_firsttransfer);
  --pio_delay_decay_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_delay_decay_s1_unreg_firsttransfer <= NOT ((pio_delay_decay_s1_slavearbiterlockenable AND pio_delay_decay_s1_any_continuerequest));
  --pio_delay_decay_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_decay_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_delay_decay_s1_begins_xfer) = '1' then 
        pio_delay_decay_s1_reg_firsttransfer <= pio_delay_decay_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_delay_decay_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_delay_decay_s1_beginbursttransfer_internal <= pio_delay_decay_s1_begins_xfer;
  --~pio_delay_decay_s1_write_n assignment, which is an e_mux
  pio_delay_decay_s1_write_n <= NOT ((((internal_cpu_data_master_granted_pio_delay_decay_s1 AND cpu_data_master_write)) AND pio_delay_decay_s1_pretend_byte_enable));
  shifted_address_to_pio_delay_decay_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_delay_decay_s1_address mux, which is an e_mux
  pio_delay_decay_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_delay_decay_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_delay_decay_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_delay_decay_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_delay_decay_s1_end_xfer <= pio_delay_decay_s1_end_xfer;
    end if;

  end process;

  --pio_delay_decay_s1_waits_for_read in a cycle, which is an e_mux
  pio_delay_decay_s1_waits_for_read <= pio_delay_decay_s1_in_a_read_cycle AND pio_delay_decay_s1_begins_xfer;
  --pio_delay_decay_s1_in_a_read_cycle assignment, which is an e_assign
  pio_delay_decay_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_delay_decay_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_delay_decay_s1_in_a_read_cycle;
  --pio_delay_decay_s1_waits_for_write in a cycle, which is an e_mux
  pio_delay_decay_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_delay_decay_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_delay_decay_s1_in_a_write_cycle assignment, which is an e_assign
  pio_delay_decay_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_delay_decay_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_delay_decay_s1_in_a_write_cycle;
  wait_for_pio_delay_decay_s1_counter <= std_logic'('0');
  --pio_delay_decay_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  pio_delay_decay_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pio_delay_decay_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_delay_decay_s1 <= internal_cpu_data_master_granted_pio_delay_decay_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_delay_decay_s1 <= internal_cpu_data_master_qualified_request_pio_delay_decay_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_delay_decay_s1 <= internal_cpu_data_master_requests_pio_delay_decay_s1;
--synthesis translate_off
    --pio_delay_decay/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_delay_length_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_delay_length_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_delay_length_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_delay_length_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_delay_length_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_delay_length_s1 : OUT STD_LOGIC;
                 signal d1_pio_delay_length_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_delay_length_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_delay_length_s1_chipselect : OUT STD_LOGIC;
                 signal pio_delay_length_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_delay_length_s1_reset_n : OUT STD_LOGIC;
                 signal pio_delay_length_s1_write_n : OUT STD_LOGIC;
                 signal pio_delay_length_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_delay_length_s1_arbitrator;


architecture europa of pio_delay_length_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_delay_length_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_delay_length_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_delay_length_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_delay_length_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_delay_length_s1 :  STD_LOGIC;
                signal pio_delay_length_s1_allgrants :  STD_LOGIC;
                signal pio_delay_length_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_delay_length_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_delay_length_s1_any_continuerequest :  STD_LOGIC;
                signal pio_delay_length_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_delay_length_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_length_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_length_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_delay_length_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_delay_length_s1_begins_xfer :  STD_LOGIC;
                signal pio_delay_length_s1_end_xfer :  STD_LOGIC;
                signal pio_delay_length_s1_firsttransfer :  STD_LOGIC;
                signal pio_delay_length_s1_grant_vector :  STD_LOGIC;
                signal pio_delay_length_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_delay_length_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_delay_length_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_delay_length_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_delay_length_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_delay_length_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_delay_length_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_delay_length_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_delay_length_s1_waits_for_read :  STD_LOGIC;
                signal pio_delay_length_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_delay_length_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_delay_length_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_delay_length_s1_end_xfer;
    end if;

  end process;

  pio_delay_length_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_delay_length_s1);
  --assign pio_delay_length_s1_readdata_from_sa = pio_delay_length_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_delay_length_s1_readdata_from_sa <= pio_delay_length_s1_readdata;
  internal_cpu_data_master_requests_pio_delay_length_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000010110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_delay_length_s1_arb_share_counter set values, which is an e_mux
  pio_delay_length_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_delay_length_s1_non_bursting_master_requests mux, which is an e_mux
  pio_delay_length_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_delay_length_s1;
  --pio_delay_length_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_delay_length_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_delay_length_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_delay_length_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_delay_length_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_delay_length_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_delay_length_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_delay_length_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_delay_length_s1_allgrants all slave grants, which is an e_mux
  pio_delay_length_s1_allgrants <= pio_delay_length_s1_grant_vector;
  --pio_delay_length_s1_end_xfer assignment, which is an e_assign
  pio_delay_length_s1_end_xfer <= NOT ((pio_delay_length_s1_waits_for_read OR pio_delay_length_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_delay_length_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_delay_length_s1 <= pio_delay_length_s1_end_xfer AND (((NOT pio_delay_length_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_delay_length_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_delay_length_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_delay_length_s1 AND pio_delay_length_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_delay_length_s1 AND NOT pio_delay_length_s1_non_bursting_master_requests));
  --pio_delay_length_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_length_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_delay_length_s1_arb_counter_enable) = '1' then 
        pio_delay_length_s1_arb_share_counter <= pio_delay_length_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_delay_length_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_length_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_delay_length_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_delay_length_s1)) OR ((end_xfer_arb_share_counter_term_pio_delay_length_s1 AND NOT pio_delay_length_s1_non_bursting_master_requests)))) = '1' then 
        pio_delay_length_s1_slavearbiterlockenable <= or_reduce(pio_delay_length_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_delay_length/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_delay_length_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_delay_length_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_delay_length_s1_slavearbiterlockenable2 <= or_reduce(pio_delay_length_s1_arb_share_counter_next_value);
  --cpu/data_master pio_delay_length/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_delay_length_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_delay_length_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_delay_length_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_delay_length_s1 <= internal_cpu_data_master_requests_pio_delay_length_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_delay_length_s1_writedata mux, which is an e_mux
  pio_delay_length_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_delay_length_s1 <= internal_cpu_data_master_qualified_request_pio_delay_length_s1;
  --cpu/data_master saved-grant pio_delay_length/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_delay_length_s1 <= internal_cpu_data_master_requests_pio_delay_length_s1;
  --allow new arb cycle for pio_delay_length/s1, which is an e_assign
  pio_delay_length_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_delay_length_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_delay_length_s1_master_qreq_vector <= std_logic'('1');
  --pio_delay_length_s1_reset_n assignment, which is an e_assign
  pio_delay_length_s1_reset_n <= reset_n;
  pio_delay_length_s1_chipselect <= internal_cpu_data_master_granted_pio_delay_length_s1;
  --pio_delay_length_s1_firsttransfer first transaction, which is an e_assign
  pio_delay_length_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_delay_length_s1_begins_xfer) = '1'), pio_delay_length_s1_unreg_firsttransfer, pio_delay_length_s1_reg_firsttransfer);
  --pio_delay_length_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_delay_length_s1_unreg_firsttransfer <= NOT ((pio_delay_length_s1_slavearbiterlockenable AND pio_delay_length_s1_any_continuerequest));
  --pio_delay_length_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_delay_length_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_delay_length_s1_begins_xfer) = '1' then 
        pio_delay_length_s1_reg_firsttransfer <= pio_delay_length_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_delay_length_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_delay_length_s1_beginbursttransfer_internal <= pio_delay_length_s1_begins_xfer;
  --~pio_delay_length_s1_write_n assignment, which is an e_mux
  pio_delay_length_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_delay_length_s1 AND cpu_data_master_write));
  shifted_address_to_pio_delay_length_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_delay_length_s1_address mux, which is an e_mux
  pio_delay_length_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_delay_length_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_delay_length_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_delay_length_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_delay_length_s1_end_xfer <= pio_delay_length_s1_end_xfer;
    end if;

  end process;

  --pio_delay_length_s1_waits_for_read in a cycle, which is an e_mux
  pio_delay_length_s1_waits_for_read <= pio_delay_length_s1_in_a_read_cycle AND pio_delay_length_s1_begins_xfer;
  --pio_delay_length_s1_in_a_read_cycle assignment, which is an e_assign
  pio_delay_length_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_delay_length_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_delay_length_s1_in_a_read_cycle;
  --pio_delay_length_s1_waits_for_write in a cycle, which is an e_mux
  pio_delay_length_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_delay_length_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_delay_length_s1_in_a_write_cycle assignment, which is an e_assign
  pio_delay_length_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_delay_length_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_delay_length_s1_in_a_write_cycle;
  wait_for_pio_delay_length_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_delay_length_s1 <= internal_cpu_data_master_granted_pio_delay_length_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_delay_length_s1 <= internal_cpu_data_master_qualified_request_pio_delay_length_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_delay_length_s1 <= internal_cpu_data_master_requests_pio_delay_length_s1;
--synthesis translate_off
    --pio_delay_length/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_master_volume_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_master_volume_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_master_volume_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_master_volume_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_master_volume_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_master_volume_s1 : OUT STD_LOGIC;
                 signal d1_pio_master_volume_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_master_volume_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_master_volume_s1_chipselect : OUT STD_LOGIC;
                 signal pio_master_volume_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_master_volume_s1_reset_n : OUT STD_LOGIC;
                 signal pio_master_volume_s1_write_n : OUT STD_LOGIC;
                 signal pio_master_volume_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_master_volume_s1_arbitrator;


architecture europa of pio_master_volume_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_master_volume_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_master_volume_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_master_volume_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_master_volume_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_master_volume_s1 :  STD_LOGIC;
                signal pio_master_volume_s1_allgrants :  STD_LOGIC;
                signal pio_master_volume_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_master_volume_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_master_volume_s1_any_continuerequest :  STD_LOGIC;
                signal pio_master_volume_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_master_volume_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_master_volume_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_master_volume_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_master_volume_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_master_volume_s1_begins_xfer :  STD_LOGIC;
                signal pio_master_volume_s1_end_xfer :  STD_LOGIC;
                signal pio_master_volume_s1_firsttransfer :  STD_LOGIC;
                signal pio_master_volume_s1_grant_vector :  STD_LOGIC;
                signal pio_master_volume_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_master_volume_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_master_volume_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_master_volume_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_master_volume_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_master_volume_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_master_volume_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_master_volume_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_master_volume_s1_waits_for_read :  STD_LOGIC;
                signal pio_master_volume_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_master_volume_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_master_volume_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_master_volume_s1_end_xfer;
    end if;

  end process;

  pio_master_volume_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_master_volume_s1);
  --assign pio_master_volume_s1_readdata_from_sa = pio_master_volume_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_master_volume_s1_readdata_from_sa <= pio_master_volume_s1_readdata;
  internal_cpu_data_master_requests_pio_master_volume_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000010100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_master_volume_s1_arb_share_counter set values, which is an e_mux
  pio_master_volume_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_master_volume_s1_non_bursting_master_requests mux, which is an e_mux
  pio_master_volume_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_master_volume_s1;
  --pio_master_volume_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_master_volume_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_master_volume_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_master_volume_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_master_volume_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_master_volume_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_master_volume_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_master_volume_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_master_volume_s1_allgrants all slave grants, which is an e_mux
  pio_master_volume_s1_allgrants <= pio_master_volume_s1_grant_vector;
  --pio_master_volume_s1_end_xfer assignment, which is an e_assign
  pio_master_volume_s1_end_xfer <= NOT ((pio_master_volume_s1_waits_for_read OR pio_master_volume_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_master_volume_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_master_volume_s1 <= pio_master_volume_s1_end_xfer AND (((NOT pio_master_volume_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_master_volume_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_master_volume_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_master_volume_s1 AND pio_master_volume_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_master_volume_s1 AND NOT pio_master_volume_s1_non_bursting_master_requests));
  --pio_master_volume_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_master_volume_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_master_volume_s1_arb_counter_enable) = '1' then 
        pio_master_volume_s1_arb_share_counter <= pio_master_volume_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_master_volume_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_master_volume_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_master_volume_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_master_volume_s1)) OR ((end_xfer_arb_share_counter_term_pio_master_volume_s1 AND NOT pio_master_volume_s1_non_bursting_master_requests)))) = '1' then 
        pio_master_volume_s1_slavearbiterlockenable <= or_reduce(pio_master_volume_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_master_volume/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_master_volume_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_master_volume_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_master_volume_s1_slavearbiterlockenable2 <= or_reduce(pio_master_volume_s1_arb_share_counter_next_value);
  --cpu/data_master pio_master_volume/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_master_volume_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_master_volume_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_master_volume_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_master_volume_s1 <= internal_cpu_data_master_requests_pio_master_volume_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_master_volume_s1_writedata mux, which is an e_mux
  pio_master_volume_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_master_volume_s1 <= internal_cpu_data_master_qualified_request_pio_master_volume_s1;
  --cpu/data_master saved-grant pio_master_volume/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_master_volume_s1 <= internal_cpu_data_master_requests_pio_master_volume_s1;
  --allow new arb cycle for pio_master_volume/s1, which is an e_assign
  pio_master_volume_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_master_volume_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_master_volume_s1_master_qreq_vector <= std_logic'('1');
  --pio_master_volume_s1_reset_n assignment, which is an e_assign
  pio_master_volume_s1_reset_n <= reset_n;
  pio_master_volume_s1_chipselect <= internal_cpu_data_master_granted_pio_master_volume_s1;
  --pio_master_volume_s1_firsttransfer first transaction, which is an e_assign
  pio_master_volume_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_master_volume_s1_begins_xfer) = '1'), pio_master_volume_s1_unreg_firsttransfer, pio_master_volume_s1_reg_firsttransfer);
  --pio_master_volume_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_master_volume_s1_unreg_firsttransfer <= NOT ((pio_master_volume_s1_slavearbiterlockenable AND pio_master_volume_s1_any_continuerequest));
  --pio_master_volume_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_master_volume_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_master_volume_s1_begins_xfer) = '1' then 
        pio_master_volume_s1_reg_firsttransfer <= pio_master_volume_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_master_volume_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_master_volume_s1_beginbursttransfer_internal <= pio_master_volume_s1_begins_xfer;
  --~pio_master_volume_s1_write_n assignment, which is an e_mux
  pio_master_volume_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_master_volume_s1 AND cpu_data_master_write));
  shifted_address_to_pio_master_volume_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_master_volume_s1_address mux, which is an e_mux
  pio_master_volume_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_master_volume_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_master_volume_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_master_volume_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_master_volume_s1_end_xfer <= pio_master_volume_s1_end_xfer;
    end if;

  end process;

  --pio_master_volume_s1_waits_for_read in a cycle, which is an e_mux
  pio_master_volume_s1_waits_for_read <= pio_master_volume_s1_in_a_read_cycle AND pio_master_volume_s1_begins_xfer;
  --pio_master_volume_s1_in_a_read_cycle assignment, which is an e_assign
  pio_master_volume_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_master_volume_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_master_volume_s1_in_a_read_cycle;
  --pio_master_volume_s1_waits_for_write in a cycle, which is an e_mux
  pio_master_volume_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_master_volume_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_master_volume_s1_in_a_write_cycle assignment, which is an e_assign
  pio_master_volume_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_master_volume_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_master_volume_s1_in_a_write_cycle;
  wait_for_pio_master_volume_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_master_volume_s1 <= internal_cpu_data_master_granted_pio_master_volume_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_master_volume_s1 <= internal_cpu_data_master_qualified_request_pio_master_volume_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_master_volume_s1 <= internal_cpu_data_master_requests_pio_master_volume_s1;
--synthesis translate_off
    --pio_master_volume/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_octaver_bypass_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_octaver_bypass_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                 signal d1_pio_octaver_bypass_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_octaver_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_octaver_bypass_s1_chipselect : OUT STD_LOGIC;
                 signal pio_octaver_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_octaver_bypass_s1_reset_n : OUT STD_LOGIC;
                 signal pio_octaver_bypass_s1_write_n : OUT STD_LOGIC;
                 signal pio_octaver_bypass_s1_writedata : OUT STD_LOGIC
              );
end entity pio_octaver_bypass_s1_arbitrator;


architecture europa of pio_octaver_bypass_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal pio_octaver_bypass_s1_allgrants :  STD_LOGIC;
                signal pio_octaver_bypass_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_octaver_bypass_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_octaver_bypass_s1_any_continuerequest :  STD_LOGIC;
                signal pio_octaver_bypass_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_octaver_bypass_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_octaver_bypass_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_octaver_bypass_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_octaver_bypass_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_octaver_bypass_s1_begins_xfer :  STD_LOGIC;
                signal pio_octaver_bypass_s1_end_xfer :  STD_LOGIC;
                signal pio_octaver_bypass_s1_firsttransfer :  STD_LOGIC;
                signal pio_octaver_bypass_s1_grant_vector :  STD_LOGIC;
                signal pio_octaver_bypass_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_octaver_bypass_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_octaver_bypass_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_octaver_bypass_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_octaver_bypass_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_octaver_bypass_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_octaver_bypass_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_octaver_bypass_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_octaver_bypass_s1_waits_for_read :  STD_LOGIC;
                signal pio_octaver_bypass_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_octaver_bypass_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_octaver_bypass_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_octaver_bypass_s1_end_xfer;
    end if;

  end process;

  pio_octaver_bypass_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_octaver_bypass_s1);
  --assign pio_octaver_bypass_s1_readdata_from_sa = pio_octaver_bypass_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_octaver_bypass_s1_readdata_from_sa <= pio_octaver_bypass_s1_readdata;
  internal_cpu_data_master_requests_pio_octaver_bypass_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000101100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_octaver_bypass_s1_arb_share_counter set values, which is an e_mux
  pio_octaver_bypass_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_octaver_bypass_s1_non_bursting_master_requests mux, which is an e_mux
  pio_octaver_bypass_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_octaver_bypass_s1;
  --pio_octaver_bypass_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_octaver_bypass_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_octaver_bypass_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_octaver_bypass_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_octaver_bypass_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_octaver_bypass_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_octaver_bypass_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_octaver_bypass_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_octaver_bypass_s1_allgrants all slave grants, which is an e_mux
  pio_octaver_bypass_s1_allgrants <= pio_octaver_bypass_s1_grant_vector;
  --pio_octaver_bypass_s1_end_xfer assignment, which is an e_assign
  pio_octaver_bypass_s1_end_xfer <= NOT ((pio_octaver_bypass_s1_waits_for_read OR pio_octaver_bypass_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_octaver_bypass_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_octaver_bypass_s1 <= pio_octaver_bypass_s1_end_xfer AND (((NOT pio_octaver_bypass_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_octaver_bypass_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_octaver_bypass_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_octaver_bypass_s1 AND pio_octaver_bypass_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_octaver_bypass_s1 AND NOT pio_octaver_bypass_s1_non_bursting_master_requests));
  --pio_octaver_bypass_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_octaver_bypass_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_octaver_bypass_s1_arb_counter_enable) = '1' then 
        pio_octaver_bypass_s1_arb_share_counter <= pio_octaver_bypass_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_octaver_bypass_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_octaver_bypass_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_octaver_bypass_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_octaver_bypass_s1)) OR ((end_xfer_arb_share_counter_term_pio_octaver_bypass_s1 AND NOT pio_octaver_bypass_s1_non_bursting_master_requests)))) = '1' then 
        pio_octaver_bypass_s1_slavearbiterlockenable <= or_reduce(pio_octaver_bypass_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_octaver_bypass/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_octaver_bypass_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_octaver_bypass_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_octaver_bypass_s1_slavearbiterlockenable2 <= or_reduce(pio_octaver_bypass_s1_arb_share_counter_next_value);
  --cpu/data_master pio_octaver_bypass/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_octaver_bypass_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_octaver_bypass_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_octaver_bypass_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_octaver_bypass_s1 <= internal_cpu_data_master_requests_pio_octaver_bypass_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_octaver_bypass_s1_writedata mux, which is an e_mux
  pio_octaver_bypass_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_octaver_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_octaver_bypass_s1;
  --cpu/data_master saved-grant pio_octaver_bypass/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_octaver_bypass_s1 <= internal_cpu_data_master_requests_pio_octaver_bypass_s1;
  --allow new arb cycle for pio_octaver_bypass/s1, which is an e_assign
  pio_octaver_bypass_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_octaver_bypass_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_octaver_bypass_s1_master_qreq_vector <= std_logic'('1');
  --pio_octaver_bypass_s1_reset_n assignment, which is an e_assign
  pio_octaver_bypass_s1_reset_n <= reset_n;
  pio_octaver_bypass_s1_chipselect <= internal_cpu_data_master_granted_pio_octaver_bypass_s1;
  --pio_octaver_bypass_s1_firsttransfer first transaction, which is an e_assign
  pio_octaver_bypass_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_octaver_bypass_s1_begins_xfer) = '1'), pio_octaver_bypass_s1_unreg_firsttransfer, pio_octaver_bypass_s1_reg_firsttransfer);
  --pio_octaver_bypass_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_octaver_bypass_s1_unreg_firsttransfer <= NOT ((pio_octaver_bypass_s1_slavearbiterlockenable AND pio_octaver_bypass_s1_any_continuerequest));
  --pio_octaver_bypass_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_octaver_bypass_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_octaver_bypass_s1_begins_xfer) = '1' then 
        pio_octaver_bypass_s1_reg_firsttransfer <= pio_octaver_bypass_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_octaver_bypass_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_octaver_bypass_s1_beginbursttransfer_internal <= pio_octaver_bypass_s1_begins_xfer;
  --~pio_octaver_bypass_s1_write_n assignment, which is an e_mux
  pio_octaver_bypass_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_octaver_bypass_s1 AND cpu_data_master_write));
  shifted_address_to_pio_octaver_bypass_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_octaver_bypass_s1_address mux, which is an e_mux
  pio_octaver_bypass_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_octaver_bypass_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_octaver_bypass_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_octaver_bypass_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_octaver_bypass_s1_end_xfer <= pio_octaver_bypass_s1_end_xfer;
    end if;

  end process;

  --pio_octaver_bypass_s1_waits_for_read in a cycle, which is an e_mux
  pio_octaver_bypass_s1_waits_for_read <= pio_octaver_bypass_s1_in_a_read_cycle AND pio_octaver_bypass_s1_begins_xfer;
  --pio_octaver_bypass_s1_in_a_read_cycle assignment, which is an e_assign
  pio_octaver_bypass_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_octaver_bypass_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_octaver_bypass_s1_in_a_read_cycle;
  --pio_octaver_bypass_s1_waits_for_write in a cycle, which is an e_mux
  pio_octaver_bypass_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_octaver_bypass_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_octaver_bypass_s1_in_a_write_cycle assignment, which is an e_assign
  pio_octaver_bypass_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_octaver_bypass_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_octaver_bypass_s1_in_a_write_cycle;
  wait_for_pio_octaver_bypass_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_octaver_bypass_s1 <= internal_cpu_data_master_granted_pio_octaver_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_octaver_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_octaver_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_octaver_bypass_s1 <= internal_cpu_data_master_requests_pio_octaver_bypass_s1;
--synthesis translate_off
    --pio_octaver_bypass/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_octaver_dry_wet_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_octaver_dry_wet_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                 signal d1_pio_octaver_dry_wet_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_octaver_dry_wet_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_octaver_dry_wet_s1_chipselect : OUT STD_LOGIC;
                 signal pio_octaver_dry_wet_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_octaver_dry_wet_s1_reset_n : OUT STD_LOGIC;
                 signal pio_octaver_dry_wet_s1_write_n : OUT STD_LOGIC;
                 signal pio_octaver_dry_wet_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_octaver_dry_wet_s1_arbitrator;


architecture europa of pio_octaver_dry_wet_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_allgrants :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_any_continuerequest :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_octaver_dry_wet_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_octaver_dry_wet_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_octaver_dry_wet_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_begins_xfer :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_end_xfer :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_firsttransfer :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_grant_vector :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_waits_for_read :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_octaver_dry_wet_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_octaver_dry_wet_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_octaver_dry_wet_s1_end_xfer;
    end if;

  end process;

  pio_octaver_dry_wet_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_octaver_dry_wet_s1);
  --assign pio_octaver_dry_wet_s1_readdata_from_sa = pio_octaver_dry_wet_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_octaver_dry_wet_s1_readdata_from_sa <= pio_octaver_dry_wet_s1_readdata;
  internal_cpu_data_master_requests_pio_octaver_dry_wet_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000101110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_octaver_dry_wet_s1_arb_share_counter set values, which is an e_mux
  pio_octaver_dry_wet_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_octaver_dry_wet_s1_non_bursting_master_requests mux, which is an e_mux
  pio_octaver_dry_wet_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_octaver_dry_wet_s1;
  --pio_octaver_dry_wet_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_octaver_dry_wet_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_octaver_dry_wet_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_octaver_dry_wet_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_octaver_dry_wet_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_octaver_dry_wet_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_octaver_dry_wet_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_octaver_dry_wet_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_octaver_dry_wet_s1_allgrants all slave grants, which is an e_mux
  pio_octaver_dry_wet_s1_allgrants <= pio_octaver_dry_wet_s1_grant_vector;
  --pio_octaver_dry_wet_s1_end_xfer assignment, which is an e_assign
  pio_octaver_dry_wet_s1_end_xfer <= NOT ((pio_octaver_dry_wet_s1_waits_for_read OR pio_octaver_dry_wet_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_octaver_dry_wet_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_octaver_dry_wet_s1 <= pio_octaver_dry_wet_s1_end_xfer AND (((NOT pio_octaver_dry_wet_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_octaver_dry_wet_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_octaver_dry_wet_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_octaver_dry_wet_s1 AND pio_octaver_dry_wet_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_octaver_dry_wet_s1 AND NOT pio_octaver_dry_wet_s1_non_bursting_master_requests));
  --pio_octaver_dry_wet_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_octaver_dry_wet_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_octaver_dry_wet_s1_arb_counter_enable) = '1' then 
        pio_octaver_dry_wet_s1_arb_share_counter <= pio_octaver_dry_wet_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_octaver_dry_wet_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_octaver_dry_wet_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_octaver_dry_wet_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_octaver_dry_wet_s1)) OR ((end_xfer_arb_share_counter_term_pio_octaver_dry_wet_s1 AND NOT pio_octaver_dry_wet_s1_non_bursting_master_requests)))) = '1' then 
        pio_octaver_dry_wet_s1_slavearbiterlockenable <= or_reduce(pio_octaver_dry_wet_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_octaver_dry_wet/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_octaver_dry_wet_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_octaver_dry_wet_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_octaver_dry_wet_s1_slavearbiterlockenable2 <= or_reduce(pio_octaver_dry_wet_s1_arb_share_counter_next_value);
  --cpu/data_master pio_octaver_dry_wet/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_octaver_dry_wet_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_octaver_dry_wet_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_octaver_dry_wet_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 <= internal_cpu_data_master_requests_pio_octaver_dry_wet_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_octaver_dry_wet_s1_writedata mux, which is an e_mux
  pio_octaver_dry_wet_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_octaver_dry_wet_s1 <= internal_cpu_data_master_qualified_request_pio_octaver_dry_wet_s1;
  --cpu/data_master saved-grant pio_octaver_dry_wet/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_octaver_dry_wet_s1 <= internal_cpu_data_master_requests_pio_octaver_dry_wet_s1;
  --allow new arb cycle for pio_octaver_dry_wet/s1, which is an e_assign
  pio_octaver_dry_wet_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_octaver_dry_wet_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_octaver_dry_wet_s1_master_qreq_vector <= std_logic'('1');
  --pio_octaver_dry_wet_s1_reset_n assignment, which is an e_assign
  pio_octaver_dry_wet_s1_reset_n <= reset_n;
  pio_octaver_dry_wet_s1_chipselect <= internal_cpu_data_master_granted_pio_octaver_dry_wet_s1;
  --pio_octaver_dry_wet_s1_firsttransfer first transaction, which is an e_assign
  pio_octaver_dry_wet_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_octaver_dry_wet_s1_begins_xfer) = '1'), pio_octaver_dry_wet_s1_unreg_firsttransfer, pio_octaver_dry_wet_s1_reg_firsttransfer);
  --pio_octaver_dry_wet_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_octaver_dry_wet_s1_unreg_firsttransfer <= NOT ((pio_octaver_dry_wet_s1_slavearbiterlockenable AND pio_octaver_dry_wet_s1_any_continuerequest));
  --pio_octaver_dry_wet_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_octaver_dry_wet_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_octaver_dry_wet_s1_begins_xfer) = '1' then 
        pio_octaver_dry_wet_s1_reg_firsttransfer <= pio_octaver_dry_wet_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_octaver_dry_wet_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_octaver_dry_wet_s1_beginbursttransfer_internal <= pio_octaver_dry_wet_s1_begins_xfer;
  --~pio_octaver_dry_wet_s1_write_n assignment, which is an e_mux
  pio_octaver_dry_wet_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_octaver_dry_wet_s1 AND cpu_data_master_write));
  shifted_address_to_pio_octaver_dry_wet_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_octaver_dry_wet_s1_address mux, which is an e_mux
  pio_octaver_dry_wet_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_octaver_dry_wet_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_octaver_dry_wet_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_octaver_dry_wet_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_octaver_dry_wet_s1_end_xfer <= pio_octaver_dry_wet_s1_end_xfer;
    end if;

  end process;

  --pio_octaver_dry_wet_s1_waits_for_read in a cycle, which is an e_mux
  pio_octaver_dry_wet_s1_waits_for_read <= pio_octaver_dry_wet_s1_in_a_read_cycle AND pio_octaver_dry_wet_s1_begins_xfer;
  --pio_octaver_dry_wet_s1_in_a_read_cycle assignment, which is an e_assign
  pio_octaver_dry_wet_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_octaver_dry_wet_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_octaver_dry_wet_s1_in_a_read_cycle;
  --pio_octaver_dry_wet_s1_waits_for_write in a cycle, which is an e_mux
  pio_octaver_dry_wet_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_octaver_dry_wet_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_octaver_dry_wet_s1_in_a_write_cycle assignment, which is an e_assign
  pio_octaver_dry_wet_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_octaver_dry_wet_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_octaver_dry_wet_s1_in_a_write_cycle;
  wait_for_pio_octaver_dry_wet_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_octaver_dry_wet_s1 <= internal_cpu_data_master_granted_pio_octaver_dry_wet_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 <= internal_cpu_data_master_qualified_request_pio_octaver_dry_wet_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_octaver_dry_wet_s1 <= internal_cpu_data_master_requests_pio_octaver_dry_wet_s1;
--synthesis translate_off
    --pio_octaver_dry_wet/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_output_power_left_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal pio_output_power_left_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_output_power_left_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_output_power_left_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_output_power_left_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_output_power_left_s1 : OUT STD_LOGIC;
                 signal d1_pio_output_power_left_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_output_power_left_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_output_power_left_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_output_power_left_s1_reset_n : OUT STD_LOGIC
              );
end entity pio_output_power_left_s1_arbitrator;


architecture europa of pio_output_power_left_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_output_power_left_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_output_power_left_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_output_power_left_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_output_power_left_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_output_power_left_s1 :  STD_LOGIC;
                signal pio_output_power_left_s1_allgrants :  STD_LOGIC;
                signal pio_output_power_left_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_output_power_left_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_output_power_left_s1_any_continuerequest :  STD_LOGIC;
                signal pio_output_power_left_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_output_power_left_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_output_power_left_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_output_power_left_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_output_power_left_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_output_power_left_s1_begins_xfer :  STD_LOGIC;
                signal pio_output_power_left_s1_end_xfer :  STD_LOGIC;
                signal pio_output_power_left_s1_firsttransfer :  STD_LOGIC;
                signal pio_output_power_left_s1_grant_vector :  STD_LOGIC;
                signal pio_output_power_left_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_output_power_left_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_output_power_left_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_output_power_left_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_output_power_left_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_output_power_left_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_output_power_left_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_output_power_left_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_output_power_left_s1_waits_for_read :  STD_LOGIC;
                signal pio_output_power_left_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_output_power_left_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_output_power_left_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_output_power_left_s1_end_xfer;
    end if;

  end process;

  pio_output_power_left_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_output_power_left_s1);
  --assign pio_output_power_left_s1_readdata_from_sa = pio_output_power_left_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_output_power_left_s1_readdata_from_sa <= pio_output_power_left_s1_readdata;
  internal_cpu_data_master_requests_pio_output_power_left_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000110000000")))) AND ((cpu_data_master_read OR cpu_data_master_write)))) AND cpu_data_master_read;
  --pio_output_power_left_s1_arb_share_counter set values, which is an e_mux
  pio_output_power_left_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_output_power_left_s1_non_bursting_master_requests mux, which is an e_mux
  pio_output_power_left_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_output_power_left_s1;
  --pio_output_power_left_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_output_power_left_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_output_power_left_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_output_power_left_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_output_power_left_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_output_power_left_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_output_power_left_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_output_power_left_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_output_power_left_s1_allgrants all slave grants, which is an e_mux
  pio_output_power_left_s1_allgrants <= pio_output_power_left_s1_grant_vector;
  --pio_output_power_left_s1_end_xfer assignment, which is an e_assign
  pio_output_power_left_s1_end_xfer <= NOT ((pio_output_power_left_s1_waits_for_read OR pio_output_power_left_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_output_power_left_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_output_power_left_s1 <= pio_output_power_left_s1_end_xfer AND (((NOT pio_output_power_left_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_output_power_left_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_output_power_left_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_output_power_left_s1 AND pio_output_power_left_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_output_power_left_s1 AND NOT pio_output_power_left_s1_non_bursting_master_requests));
  --pio_output_power_left_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_output_power_left_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_output_power_left_s1_arb_counter_enable) = '1' then 
        pio_output_power_left_s1_arb_share_counter <= pio_output_power_left_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_output_power_left_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_output_power_left_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_output_power_left_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_output_power_left_s1)) OR ((end_xfer_arb_share_counter_term_pio_output_power_left_s1 AND NOT pio_output_power_left_s1_non_bursting_master_requests)))) = '1' then 
        pio_output_power_left_s1_slavearbiterlockenable <= or_reduce(pio_output_power_left_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_output_power_left/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_output_power_left_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_output_power_left_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_output_power_left_s1_slavearbiterlockenable2 <= or_reduce(pio_output_power_left_s1_arb_share_counter_next_value);
  --cpu/data_master pio_output_power_left/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_output_power_left_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_output_power_left_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_output_power_left_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_output_power_left_s1 <= internal_cpu_data_master_requests_pio_output_power_left_s1;
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_output_power_left_s1 <= internal_cpu_data_master_qualified_request_pio_output_power_left_s1;
  --cpu/data_master saved-grant pio_output_power_left/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_output_power_left_s1 <= internal_cpu_data_master_requests_pio_output_power_left_s1;
  --allow new arb cycle for pio_output_power_left/s1, which is an e_assign
  pio_output_power_left_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_output_power_left_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_output_power_left_s1_master_qreq_vector <= std_logic'('1');
  --pio_output_power_left_s1_reset_n assignment, which is an e_assign
  pio_output_power_left_s1_reset_n <= reset_n;
  --pio_output_power_left_s1_firsttransfer first transaction, which is an e_assign
  pio_output_power_left_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_output_power_left_s1_begins_xfer) = '1'), pio_output_power_left_s1_unreg_firsttransfer, pio_output_power_left_s1_reg_firsttransfer);
  --pio_output_power_left_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_output_power_left_s1_unreg_firsttransfer <= NOT ((pio_output_power_left_s1_slavearbiterlockenable AND pio_output_power_left_s1_any_continuerequest));
  --pio_output_power_left_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_output_power_left_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_output_power_left_s1_begins_xfer) = '1' then 
        pio_output_power_left_s1_reg_firsttransfer <= pio_output_power_left_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_output_power_left_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_output_power_left_s1_beginbursttransfer_internal <= pio_output_power_left_s1_begins_xfer;
  shifted_address_to_pio_output_power_left_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_output_power_left_s1_address mux, which is an e_mux
  pio_output_power_left_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_output_power_left_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_output_power_left_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_output_power_left_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_output_power_left_s1_end_xfer <= pio_output_power_left_s1_end_xfer;
    end if;

  end process;

  --pio_output_power_left_s1_waits_for_read in a cycle, which is an e_mux
  pio_output_power_left_s1_waits_for_read <= pio_output_power_left_s1_in_a_read_cycle AND pio_output_power_left_s1_begins_xfer;
  --pio_output_power_left_s1_in_a_read_cycle assignment, which is an e_assign
  pio_output_power_left_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_output_power_left_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_output_power_left_s1_in_a_read_cycle;
  --pio_output_power_left_s1_waits_for_write in a cycle, which is an e_mux
  pio_output_power_left_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_output_power_left_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_output_power_left_s1_in_a_write_cycle assignment, which is an e_assign
  pio_output_power_left_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_output_power_left_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_output_power_left_s1_in_a_write_cycle;
  wait_for_pio_output_power_left_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_output_power_left_s1 <= internal_cpu_data_master_granted_pio_output_power_left_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_output_power_left_s1 <= internal_cpu_data_master_qualified_request_pio_output_power_left_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_output_power_left_s1 <= internal_cpu_data_master_requests_pio_output_power_left_s1;
--synthesis translate_off
    --pio_output_power_left/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_output_power_right_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal pio_output_power_right_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_output_power_right_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_output_power_right_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_output_power_right_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_output_power_right_s1 : OUT STD_LOGIC;
                 signal d1_pio_output_power_right_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_output_power_right_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_output_power_right_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_output_power_right_s1_reset_n : OUT STD_LOGIC
              );
end entity pio_output_power_right_s1_arbitrator;


architecture europa of pio_output_power_right_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_output_power_right_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_output_power_right_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_output_power_right_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_output_power_right_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_output_power_right_s1 :  STD_LOGIC;
                signal pio_output_power_right_s1_allgrants :  STD_LOGIC;
                signal pio_output_power_right_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_output_power_right_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_output_power_right_s1_any_continuerequest :  STD_LOGIC;
                signal pio_output_power_right_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_output_power_right_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_output_power_right_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_output_power_right_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_output_power_right_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_output_power_right_s1_begins_xfer :  STD_LOGIC;
                signal pio_output_power_right_s1_end_xfer :  STD_LOGIC;
                signal pio_output_power_right_s1_firsttransfer :  STD_LOGIC;
                signal pio_output_power_right_s1_grant_vector :  STD_LOGIC;
                signal pio_output_power_right_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_output_power_right_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_output_power_right_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_output_power_right_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_output_power_right_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_output_power_right_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_output_power_right_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_output_power_right_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_output_power_right_s1_waits_for_read :  STD_LOGIC;
                signal pio_output_power_right_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_output_power_right_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_output_power_right_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_output_power_right_s1_end_xfer;
    end if;

  end process;

  pio_output_power_right_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_output_power_right_s1);
  --assign pio_output_power_right_s1_readdata_from_sa = pio_output_power_right_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_output_power_right_s1_readdata_from_sa <= pio_output_power_right_s1_readdata;
  internal_cpu_data_master_requests_pio_output_power_right_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000110100000")))) AND ((cpu_data_master_read OR cpu_data_master_write)))) AND cpu_data_master_read;
  --pio_output_power_right_s1_arb_share_counter set values, which is an e_mux
  pio_output_power_right_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_output_power_right_s1_non_bursting_master_requests mux, which is an e_mux
  pio_output_power_right_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_output_power_right_s1;
  --pio_output_power_right_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_output_power_right_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_output_power_right_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_output_power_right_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_output_power_right_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_output_power_right_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_output_power_right_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_output_power_right_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_output_power_right_s1_allgrants all slave grants, which is an e_mux
  pio_output_power_right_s1_allgrants <= pio_output_power_right_s1_grant_vector;
  --pio_output_power_right_s1_end_xfer assignment, which is an e_assign
  pio_output_power_right_s1_end_xfer <= NOT ((pio_output_power_right_s1_waits_for_read OR pio_output_power_right_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_output_power_right_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_output_power_right_s1 <= pio_output_power_right_s1_end_xfer AND (((NOT pio_output_power_right_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_output_power_right_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_output_power_right_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_output_power_right_s1 AND pio_output_power_right_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_output_power_right_s1 AND NOT pio_output_power_right_s1_non_bursting_master_requests));
  --pio_output_power_right_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_output_power_right_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_output_power_right_s1_arb_counter_enable) = '1' then 
        pio_output_power_right_s1_arb_share_counter <= pio_output_power_right_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_output_power_right_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_output_power_right_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_output_power_right_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_output_power_right_s1)) OR ((end_xfer_arb_share_counter_term_pio_output_power_right_s1 AND NOT pio_output_power_right_s1_non_bursting_master_requests)))) = '1' then 
        pio_output_power_right_s1_slavearbiterlockenable <= or_reduce(pio_output_power_right_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_output_power_right/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_output_power_right_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_output_power_right_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_output_power_right_s1_slavearbiterlockenable2 <= or_reduce(pio_output_power_right_s1_arb_share_counter_next_value);
  --cpu/data_master pio_output_power_right/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_output_power_right_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_output_power_right_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_output_power_right_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_output_power_right_s1 <= internal_cpu_data_master_requests_pio_output_power_right_s1;
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_output_power_right_s1 <= internal_cpu_data_master_qualified_request_pio_output_power_right_s1;
  --cpu/data_master saved-grant pio_output_power_right/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_output_power_right_s1 <= internal_cpu_data_master_requests_pio_output_power_right_s1;
  --allow new arb cycle for pio_output_power_right/s1, which is an e_assign
  pio_output_power_right_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_output_power_right_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_output_power_right_s1_master_qreq_vector <= std_logic'('1');
  --pio_output_power_right_s1_reset_n assignment, which is an e_assign
  pio_output_power_right_s1_reset_n <= reset_n;
  --pio_output_power_right_s1_firsttransfer first transaction, which is an e_assign
  pio_output_power_right_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_output_power_right_s1_begins_xfer) = '1'), pio_output_power_right_s1_unreg_firsttransfer, pio_output_power_right_s1_reg_firsttransfer);
  --pio_output_power_right_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_output_power_right_s1_unreg_firsttransfer <= NOT ((pio_output_power_right_s1_slavearbiterlockenable AND pio_output_power_right_s1_any_continuerequest));
  --pio_output_power_right_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_output_power_right_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_output_power_right_s1_begins_xfer) = '1' then 
        pio_output_power_right_s1_reg_firsttransfer <= pio_output_power_right_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_output_power_right_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_output_power_right_s1_beginbursttransfer_internal <= pio_output_power_right_s1_begins_xfer;
  shifted_address_to_pio_output_power_right_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_output_power_right_s1_address mux, which is an e_mux
  pio_output_power_right_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_output_power_right_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_output_power_right_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_output_power_right_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_output_power_right_s1_end_xfer <= pio_output_power_right_s1_end_xfer;
    end if;

  end process;

  --pio_output_power_right_s1_waits_for_read in a cycle, which is an e_mux
  pio_output_power_right_s1_waits_for_read <= pio_output_power_right_s1_in_a_read_cycle AND pio_output_power_right_s1_begins_xfer;
  --pio_output_power_right_s1_in_a_read_cycle assignment, which is an e_assign
  pio_output_power_right_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_output_power_right_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_output_power_right_s1_in_a_read_cycle;
  --pio_output_power_right_s1_waits_for_write in a cycle, which is an e_mux
  pio_output_power_right_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_output_power_right_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_output_power_right_s1_in_a_write_cycle assignment, which is an e_assign
  pio_output_power_right_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_output_power_right_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_output_power_right_s1_in_a_write_cycle;
  wait_for_pio_output_power_right_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_output_power_right_s1 <= internal_cpu_data_master_granted_pio_output_power_right_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_output_power_right_s1 <= internal_cpu_data_master_qualified_request_pio_output_power_right_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_output_power_right_s1 <= internal_cpu_data_master_requests_pio_output_power_right_s1;
--synthesis translate_off
    --pio_output_power_right/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_overdrive_asymmetric_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_overdrive_asymmetric_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                 signal d1_pio_overdrive_asymmetric_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_overdrive_asymmetric_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_overdrive_asymmetric_s1_chipselect : OUT STD_LOGIC;
                 signal pio_overdrive_asymmetric_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_overdrive_asymmetric_s1_reset_n : OUT STD_LOGIC;
                 signal pio_overdrive_asymmetric_s1_write_n : OUT STD_LOGIC;
                 signal pio_overdrive_asymmetric_s1_writedata : OUT STD_LOGIC
              );
end entity pio_overdrive_asymmetric_s1_arbitrator;


architecture europa of pio_overdrive_asymmetric_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_allgrants :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_any_continuerequest :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_asymmetric_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_asymmetric_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_asymmetric_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_begins_xfer :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_end_xfer :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_grant_vector :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_waits_for_read :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_overdrive_asymmetric_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_overdrive_asymmetric_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_overdrive_asymmetric_s1_end_xfer;
    end if;

  end process;

  pio_overdrive_asymmetric_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1);
  --assign pio_overdrive_asymmetric_s1_readdata_from_sa = pio_overdrive_asymmetric_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_overdrive_asymmetric_s1_readdata_from_sa <= pio_overdrive_asymmetric_s1_readdata;
  internal_cpu_data_master_requests_pio_overdrive_asymmetric_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000001110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_overdrive_asymmetric_s1_arb_share_counter set values, which is an e_mux
  pio_overdrive_asymmetric_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_overdrive_asymmetric_s1_non_bursting_master_requests mux, which is an e_mux
  pio_overdrive_asymmetric_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_overdrive_asymmetric_s1;
  --pio_overdrive_asymmetric_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_overdrive_asymmetric_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_overdrive_asymmetric_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_overdrive_asymmetric_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_overdrive_asymmetric_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_asymmetric_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_overdrive_asymmetric_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_asymmetric_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_overdrive_asymmetric_s1_allgrants all slave grants, which is an e_mux
  pio_overdrive_asymmetric_s1_allgrants <= pio_overdrive_asymmetric_s1_grant_vector;
  --pio_overdrive_asymmetric_s1_end_xfer assignment, which is an e_assign
  pio_overdrive_asymmetric_s1_end_xfer <= NOT ((pio_overdrive_asymmetric_s1_waits_for_read OR pio_overdrive_asymmetric_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_overdrive_asymmetric_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_overdrive_asymmetric_s1 <= pio_overdrive_asymmetric_s1_end_xfer AND (((NOT pio_overdrive_asymmetric_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_overdrive_asymmetric_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_overdrive_asymmetric_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_overdrive_asymmetric_s1 AND pio_overdrive_asymmetric_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_asymmetric_s1 AND NOT pio_overdrive_asymmetric_s1_non_bursting_master_requests));
  --pio_overdrive_asymmetric_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_asymmetric_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_asymmetric_s1_arb_counter_enable) = '1' then 
        pio_overdrive_asymmetric_s1_arb_share_counter <= pio_overdrive_asymmetric_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_overdrive_asymmetric_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_asymmetric_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_overdrive_asymmetric_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_overdrive_asymmetric_s1)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_asymmetric_s1 AND NOT pio_overdrive_asymmetric_s1_non_bursting_master_requests)))) = '1' then 
        pio_overdrive_asymmetric_s1_slavearbiterlockenable <= or_reduce(pio_overdrive_asymmetric_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_overdrive_asymmetric/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_overdrive_asymmetric_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_overdrive_asymmetric_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_overdrive_asymmetric_s1_slavearbiterlockenable2 <= or_reduce(pio_overdrive_asymmetric_s1_arb_share_counter_next_value);
  --cpu/data_master pio_overdrive_asymmetric/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_overdrive_asymmetric_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_overdrive_asymmetric_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_overdrive_asymmetric_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 <= internal_cpu_data_master_requests_pio_overdrive_asymmetric_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_overdrive_asymmetric_s1_writedata mux, which is an e_mux
  pio_overdrive_asymmetric_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_overdrive_asymmetric_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1;
  --cpu/data_master saved-grant pio_overdrive_asymmetric/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_overdrive_asymmetric_s1 <= internal_cpu_data_master_requests_pio_overdrive_asymmetric_s1;
  --allow new arb cycle for pio_overdrive_asymmetric/s1, which is an e_assign
  pio_overdrive_asymmetric_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_overdrive_asymmetric_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_overdrive_asymmetric_s1_master_qreq_vector <= std_logic'('1');
  --pio_overdrive_asymmetric_s1_reset_n assignment, which is an e_assign
  pio_overdrive_asymmetric_s1_reset_n <= reset_n;
  pio_overdrive_asymmetric_s1_chipselect <= internal_cpu_data_master_granted_pio_overdrive_asymmetric_s1;
  --pio_overdrive_asymmetric_s1_firsttransfer first transaction, which is an e_assign
  pio_overdrive_asymmetric_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_overdrive_asymmetric_s1_begins_xfer) = '1'), pio_overdrive_asymmetric_s1_unreg_firsttransfer, pio_overdrive_asymmetric_s1_reg_firsttransfer);
  --pio_overdrive_asymmetric_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_overdrive_asymmetric_s1_unreg_firsttransfer <= NOT ((pio_overdrive_asymmetric_s1_slavearbiterlockenable AND pio_overdrive_asymmetric_s1_any_continuerequest));
  --pio_overdrive_asymmetric_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_asymmetric_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_asymmetric_s1_begins_xfer) = '1' then 
        pio_overdrive_asymmetric_s1_reg_firsttransfer <= pio_overdrive_asymmetric_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_overdrive_asymmetric_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_overdrive_asymmetric_s1_beginbursttransfer_internal <= pio_overdrive_asymmetric_s1_begins_xfer;
  --~pio_overdrive_asymmetric_s1_write_n assignment, which is an e_mux
  pio_overdrive_asymmetric_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_overdrive_asymmetric_s1 AND cpu_data_master_write));
  shifted_address_to_pio_overdrive_asymmetric_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_overdrive_asymmetric_s1_address mux, which is an e_mux
  pio_overdrive_asymmetric_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_overdrive_asymmetric_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_overdrive_asymmetric_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_overdrive_asymmetric_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_overdrive_asymmetric_s1_end_xfer <= pio_overdrive_asymmetric_s1_end_xfer;
    end if;

  end process;

  --pio_overdrive_asymmetric_s1_waits_for_read in a cycle, which is an e_mux
  pio_overdrive_asymmetric_s1_waits_for_read <= pio_overdrive_asymmetric_s1_in_a_read_cycle AND pio_overdrive_asymmetric_s1_begins_xfer;
  --pio_overdrive_asymmetric_s1_in_a_read_cycle assignment, which is an e_assign
  pio_overdrive_asymmetric_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_overdrive_asymmetric_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_overdrive_asymmetric_s1_in_a_read_cycle;
  --pio_overdrive_asymmetric_s1_waits_for_write in a cycle, which is an e_mux
  pio_overdrive_asymmetric_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_overdrive_asymmetric_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_overdrive_asymmetric_s1_in_a_write_cycle assignment, which is an e_assign
  pio_overdrive_asymmetric_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_overdrive_asymmetric_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_overdrive_asymmetric_s1_in_a_write_cycle;
  wait_for_pio_overdrive_asymmetric_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_overdrive_asymmetric_s1 <= internal_cpu_data_master_granted_pio_overdrive_asymmetric_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_overdrive_asymmetric_s1 <= internal_cpu_data_master_requests_pio_overdrive_asymmetric_s1;
--synthesis translate_off
    --pio_overdrive_asymmetric/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_overdrive_bypass_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_overdrive_bypass_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                 signal d1_pio_overdrive_bypass_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_overdrive_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_overdrive_bypass_s1_chipselect : OUT STD_LOGIC;
                 signal pio_overdrive_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_overdrive_bypass_s1_reset_n : OUT STD_LOGIC;
                 signal pio_overdrive_bypass_s1_write_n : OUT STD_LOGIC;
                 signal pio_overdrive_bypass_s1_writedata : OUT STD_LOGIC
              );
end entity pio_overdrive_bypass_s1_arbitrator;


architecture europa of pio_overdrive_bypass_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_allgrants :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_any_continuerequest :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_bypass_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_bypass_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_bypass_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_begins_xfer :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_end_xfer :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_grant_vector :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_waits_for_read :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_overdrive_bypass_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_overdrive_bypass_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_overdrive_bypass_s1_end_xfer;
    end if;

  end process;

  pio_overdrive_bypass_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_overdrive_bypass_s1);
  --assign pio_overdrive_bypass_s1_readdata_from_sa = pio_overdrive_bypass_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_overdrive_bypass_s1_readdata_from_sa <= pio_overdrive_bypass_s1_readdata;
  internal_cpu_data_master_requests_pio_overdrive_bypass_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000001100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_overdrive_bypass_s1_arb_share_counter set values, which is an e_mux
  pio_overdrive_bypass_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_overdrive_bypass_s1_non_bursting_master_requests mux, which is an e_mux
  pio_overdrive_bypass_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_overdrive_bypass_s1;
  --pio_overdrive_bypass_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_overdrive_bypass_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_overdrive_bypass_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_overdrive_bypass_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_overdrive_bypass_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_bypass_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_overdrive_bypass_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_bypass_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_overdrive_bypass_s1_allgrants all slave grants, which is an e_mux
  pio_overdrive_bypass_s1_allgrants <= pio_overdrive_bypass_s1_grant_vector;
  --pio_overdrive_bypass_s1_end_xfer assignment, which is an e_assign
  pio_overdrive_bypass_s1_end_xfer <= NOT ((pio_overdrive_bypass_s1_waits_for_read OR pio_overdrive_bypass_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_overdrive_bypass_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_overdrive_bypass_s1 <= pio_overdrive_bypass_s1_end_xfer AND (((NOT pio_overdrive_bypass_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_overdrive_bypass_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_overdrive_bypass_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_overdrive_bypass_s1 AND pio_overdrive_bypass_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_bypass_s1 AND NOT pio_overdrive_bypass_s1_non_bursting_master_requests));
  --pio_overdrive_bypass_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_bypass_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_bypass_s1_arb_counter_enable) = '1' then 
        pio_overdrive_bypass_s1_arb_share_counter <= pio_overdrive_bypass_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_overdrive_bypass_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_bypass_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_overdrive_bypass_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_overdrive_bypass_s1)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_bypass_s1 AND NOT pio_overdrive_bypass_s1_non_bursting_master_requests)))) = '1' then 
        pio_overdrive_bypass_s1_slavearbiterlockenable <= or_reduce(pio_overdrive_bypass_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_overdrive_bypass/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_overdrive_bypass_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_overdrive_bypass_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_overdrive_bypass_s1_slavearbiterlockenable2 <= or_reduce(pio_overdrive_bypass_s1_arb_share_counter_next_value);
  --cpu/data_master pio_overdrive_bypass/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_overdrive_bypass_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_overdrive_bypass_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_overdrive_bypass_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_overdrive_bypass_s1 <= internal_cpu_data_master_requests_pio_overdrive_bypass_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_overdrive_bypass_s1_writedata mux, which is an e_mux
  pio_overdrive_bypass_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_overdrive_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_bypass_s1;
  --cpu/data_master saved-grant pio_overdrive_bypass/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_overdrive_bypass_s1 <= internal_cpu_data_master_requests_pio_overdrive_bypass_s1;
  --allow new arb cycle for pio_overdrive_bypass/s1, which is an e_assign
  pio_overdrive_bypass_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_overdrive_bypass_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_overdrive_bypass_s1_master_qreq_vector <= std_logic'('1');
  --pio_overdrive_bypass_s1_reset_n assignment, which is an e_assign
  pio_overdrive_bypass_s1_reset_n <= reset_n;
  pio_overdrive_bypass_s1_chipselect <= internal_cpu_data_master_granted_pio_overdrive_bypass_s1;
  --pio_overdrive_bypass_s1_firsttransfer first transaction, which is an e_assign
  pio_overdrive_bypass_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_overdrive_bypass_s1_begins_xfer) = '1'), pio_overdrive_bypass_s1_unreg_firsttransfer, pio_overdrive_bypass_s1_reg_firsttransfer);
  --pio_overdrive_bypass_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_overdrive_bypass_s1_unreg_firsttransfer <= NOT ((pio_overdrive_bypass_s1_slavearbiterlockenable AND pio_overdrive_bypass_s1_any_continuerequest));
  --pio_overdrive_bypass_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_bypass_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_bypass_s1_begins_xfer) = '1' then 
        pio_overdrive_bypass_s1_reg_firsttransfer <= pio_overdrive_bypass_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_overdrive_bypass_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_overdrive_bypass_s1_beginbursttransfer_internal <= pio_overdrive_bypass_s1_begins_xfer;
  --~pio_overdrive_bypass_s1_write_n assignment, which is an e_mux
  pio_overdrive_bypass_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_overdrive_bypass_s1 AND cpu_data_master_write));
  shifted_address_to_pio_overdrive_bypass_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_overdrive_bypass_s1_address mux, which is an e_mux
  pio_overdrive_bypass_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_overdrive_bypass_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_overdrive_bypass_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_overdrive_bypass_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_overdrive_bypass_s1_end_xfer <= pio_overdrive_bypass_s1_end_xfer;
    end if;

  end process;

  --pio_overdrive_bypass_s1_waits_for_read in a cycle, which is an e_mux
  pio_overdrive_bypass_s1_waits_for_read <= pio_overdrive_bypass_s1_in_a_read_cycle AND pio_overdrive_bypass_s1_begins_xfer;
  --pio_overdrive_bypass_s1_in_a_read_cycle assignment, which is an e_assign
  pio_overdrive_bypass_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_overdrive_bypass_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_overdrive_bypass_s1_in_a_read_cycle;
  --pio_overdrive_bypass_s1_waits_for_write in a cycle, which is an e_mux
  pio_overdrive_bypass_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_overdrive_bypass_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_overdrive_bypass_s1_in_a_write_cycle assignment, which is an e_assign
  pio_overdrive_bypass_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_overdrive_bypass_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_overdrive_bypass_s1_in_a_write_cycle;
  wait_for_pio_overdrive_bypass_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_overdrive_bypass_s1 <= internal_cpu_data_master_granted_pio_overdrive_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_overdrive_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_overdrive_bypass_s1 <= internal_cpu_data_master_requests_pio_overdrive_bypass_s1;
--synthesis translate_off
    --pio_overdrive_bypass/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_overdrive_gain_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_overdrive_gain_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                 signal d1_pio_overdrive_gain_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_overdrive_gain_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_overdrive_gain_s1_chipselect : OUT STD_LOGIC;
                 signal pio_overdrive_gain_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_overdrive_gain_s1_reset_n : OUT STD_LOGIC;
                 signal pio_overdrive_gain_s1_write_n : OUT STD_LOGIC;
                 signal pio_overdrive_gain_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_overdrive_gain_s1_arbitrator;


architecture europa of pio_overdrive_gain_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal pio_overdrive_gain_s1_allgrants :  STD_LOGIC;
                signal pio_overdrive_gain_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_overdrive_gain_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_overdrive_gain_s1_any_continuerequest :  STD_LOGIC;
                signal pio_overdrive_gain_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_overdrive_gain_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_gain_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_gain_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_gain_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_overdrive_gain_s1_begins_xfer :  STD_LOGIC;
                signal pio_overdrive_gain_s1_end_xfer :  STD_LOGIC;
                signal pio_overdrive_gain_s1_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_gain_s1_grant_vector :  STD_LOGIC;
                signal pio_overdrive_gain_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_overdrive_gain_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_overdrive_gain_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_overdrive_gain_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_overdrive_gain_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_gain_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_overdrive_gain_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_overdrive_gain_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_gain_s1_waits_for_read :  STD_LOGIC;
                signal pio_overdrive_gain_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_overdrive_gain_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_overdrive_gain_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_overdrive_gain_s1_end_xfer;
    end if;

  end process;

  pio_overdrive_gain_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_overdrive_gain_s1);
  --assign pio_overdrive_gain_s1_readdata_from_sa = pio_overdrive_gain_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_overdrive_gain_s1_readdata_from_sa <= pio_overdrive_gain_s1_readdata;
  internal_cpu_data_master_requests_pio_overdrive_gain_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000010010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_overdrive_gain_s1_arb_share_counter set values, which is an e_mux
  pio_overdrive_gain_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_overdrive_gain_s1_non_bursting_master_requests mux, which is an e_mux
  pio_overdrive_gain_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_overdrive_gain_s1;
  --pio_overdrive_gain_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_overdrive_gain_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_overdrive_gain_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_overdrive_gain_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_overdrive_gain_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_gain_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_overdrive_gain_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_gain_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_overdrive_gain_s1_allgrants all slave grants, which is an e_mux
  pio_overdrive_gain_s1_allgrants <= pio_overdrive_gain_s1_grant_vector;
  --pio_overdrive_gain_s1_end_xfer assignment, which is an e_assign
  pio_overdrive_gain_s1_end_xfer <= NOT ((pio_overdrive_gain_s1_waits_for_read OR pio_overdrive_gain_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_overdrive_gain_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_overdrive_gain_s1 <= pio_overdrive_gain_s1_end_xfer AND (((NOT pio_overdrive_gain_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_overdrive_gain_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_overdrive_gain_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_overdrive_gain_s1 AND pio_overdrive_gain_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_gain_s1 AND NOT pio_overdrive_gain_s1_non_bursting_master_requests));
  --pio_overdrive_gain_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_gain_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_gain_s1_arb_counter_enable) = '1' then 
        pio_overdrive_gain_s1_arb_share_counter <= pio_overdrive_gain_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_overdrive_gain_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_gain_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_overdrive_gain_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_overdrive_gain_s1)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_gain_s1 AND NOT pio_overdrive_gain_s1_non_bursting_master_requests)))) = '1' then 
        pio_overdrive_gain_s1_slavearbiterlockenable <= or_reduce(pio_overdrive_gain_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_overdrive_gain/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_overdrive_gain_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_overdrive_gain_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_overdrive_gain_s1_slavearbiterlockenable2 <= or_reduce(pio_overdrive_gain_s1_arb_share_counter_next_value);
  --cpu/data_master pio_overdrive_gain/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_overdrive_gain_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_overdrive_gain_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_overdrive_gain_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_overdrive_gain_s1 <= internal_cpu_data_master_requests_pio_overdrive_gain_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_overdrive_gain_s1_writedata mux, which is an e_mux
  pio_overdrive_gain_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_overdrive_gain_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_gain_s1;
  --cpu/data_master saved-grant pio_overdrive_gain/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_overdrive_gain_s1 <= internal_cpu_data_master_requests_pio_overdrive_gain_s1;
  --allow new arb cycle for pio_overdrive_gain/s1, which is an e_assign
  pio_overdrive_gain_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_overdrive_gain_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_overdrive_gain_s1_master_qreq_vector <= std_logic'('1');
  --pio_overdrive_gain_s1_reset_n assignment, which is an e_assign
  pio_overdrive_gain_s1_reset_n <= reset_n;
  pio_overdrive_gain_s1_chipselect <= internal_cpu_data_master_granted_pio_overdrive_gain_s1;
  --pio_overdrive_gain_s1_firsttransfer first transaction, which is an e_assign
  pio_overdrive_gain_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_overdrive_gain_s1_begins_xfer) = '1'), pio_overdrive_gain_s1_unreg_firsttransfer, pio_overdrive_gain_s1_reg_firsttransfer);
  --pio_overdrive_gain_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_overdrive_gain_s1_unreg_firsttransfer <= NOT ((pio_overdrive_gain_s1_slavearbiterlockenable AND pio_overdrive_gain_s1_any_continuerequest));
  --pio_overdrive_gain_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_gain_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_gain_s1_begins_xfer) = '1' then 
        pio_overdrive_gain_s1_reg_firsttransfer <= pio_overdrive_gain_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_overdrive_gain_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_overdrive_gain_s1_beginbursttransfer_internal <= pio_overdrive_gain_s1_begins_xfer;
  --~pio_overdrive_gain_s1_write_n assignment, which is an e_mux
  pio_overdrive_gain_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_overdrive_gain_s1 AND cpu_data_master_write));
  shifted_address_to_pio_overdrive_gain_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_overdrive_gain_s1_address mux, which is an e_mux
  pio_overdrive_gain_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_overdrive_gain_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_overdrive_gain_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_overdrive_gain_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_overdrive_gain_s1_end_xfer <= pio_overdrive_gain_s1_end_xfer;
    end if;

  end process;

  --pio_overdrive_gain_s1_waits_for_read in a cycle, which is an e_mux
  pio_overdrive_gain_s1_waits_for_read <= pio_overdrive_gain_s1_in_a_read_cycle AND pio_overdrive_gain_s1_begins_xfer;
  --pio_overdrive_gain_s1_in_a_read_cycle assignment, which is an e_assign
  pio_overdrive_gain_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_overdrive_gain_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_overdrive_gain_s1_in_a_read_cycle;
  --pio_overdrive_gain_s1_waits_for_write in a cycle, which is an e_mux
  pio_overdrive_gain_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_overdrive_gain_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_overdrive_gain_s1_in_a_write_cycle assignment, which is an e_assign
  pio_overdrive_gain_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_overdrive_gain_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_overdrive_gain_s1_in_a_write_cycle;
  wait_for_pio_overdrive_gain_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_overdrive_gain_s1 <= internal_cpu_data_master_granted_pio_overdrive_gain_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_overdrive_gain_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_gain_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_overdrive_gain_s1 <= internal_cpu_data_master_requests_pio_overdrive_gain_s1;
--synthesis translate_off
    --pio_overdrive_gain/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_overdrive_tone_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_overdrive_tone_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                 signal d1_pio_overdrive_tone_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_overdrive_tone_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_overdrive_tone_s1_chipselect : OUT STD_LOGIC;
                 signal pio_overdrive_tone_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_overdrive_tone_s1_reset_n : OUT STD_LOGIC;
                 signal pio_overdrive_tone_s1_write_n : OUT STD_LOGIC;
                 signal pio_overdrive_tone_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_overdrive_tone_s1_arbitrator;


architecture europa of pio_overdrive_tone_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal pio_overdrive_tone_s1_allgrants :  STD_LOGIC;
                signal pio_overdrive_tone_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_overdrive_tone_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_overdrive_tone_s1_any_continuerequest :  STD_LOGIC;
                signal pio_overdrive_tone_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_overdrive_tone_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_tone_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_tone_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_tone_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_overdrive_tone_s1_begins_xfer :  STD_LOGIC;
                signal pio_overdrive_tone_s1_end_xfer :  STD_LOGIC;
                signal pio_overdrive_tone_s1_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_tone_s1_grant_vector :  STD_LOGIC;
                signal pio_overdrive_tone_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_overdrive_tone_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_overdrive_tone_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_overdrive_tone_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_overdrive_tone_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_tone_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_overdrive_tone_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_overdrive_tone_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_tone_s1_waits_for_read :  STD_LOGIC;
                signal pio_overdrive_tone_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_overdrive_tone_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_overdrive_tone_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_overdrive_tone_s1_end_xfer;
    end if;

  end process;

  pio_overdrive_tone_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_overdrive_tone_s1);
  --assign pio_overdrive_tone_s1_readdata_from_sa = pio_overdrive_tone_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_overdrive_tone_s1_readdata_from_sa <= pio_overdrive_tone_s1_readdata;
  internal_cpu_data_master_requests_pio_overdrive_tone_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000001000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_overdrive_tone_s1_arb_share_counter set values, which is an e_mux
  pio_overdrive_tone_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_overdrive_tone_s1_non_bursting_master_requests mux, which is an e_mux
  pio_overdrive_tone_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_overdrive_tone_s1;
  --pio_overdrive_tone_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_overdrive_tone_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_overdrive_tone_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_overdrive_tone_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_overdrive_tone_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_tone_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_overdrive_tone_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_tone_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_overdrive_tone_s1_allgrants all slave grants, which is an e_mux
  pio_overdrive_tone_s1_allgrants <= pio_overdrive_tone_s1_grant_vector;
  --pio_overdrive_tone_s1_end_xfer assignment, which is an e_assign
  pio_overdrive_tone_s1_end_xfer <= NOT ((pio_overdrive_tone_s1_waits_for_read OR pio_overdrive_tone_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_overdrive_tone_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_overdrive_tone_s1 <= pio_overdrive_tone_s1_end_xfer AND (((NOT pio_overdrive_tone_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_overdrive_tone_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_overdrive_tone_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_overdrive_tone_s1 AND pio_overdrive_tone_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_tone_s1 AND NOT pio_overdrive_tone_s1_non_bursting_master_requests));
  --pio_overdrive_tone_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_tone_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_tone_s1_arb_counter_enable) = '1' then 
        pio_overdrive_tone_s1_arb_share_counter <= pio_overdrive_tone_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_overdrive_tone_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_tone_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_overdrive_tone_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_overdrive_tone_s1)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_tone_s1 AND NOT pio_overdrive_tone_s1_non_bursting_master_requests)))) = '1' then 
        pio_overdrive_tone_s1_slavearbiterlockenable <= or_reduce(pio_overdrive_tone_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_overdrive_tone/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_overdrive_tone_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_overdrive_tone_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_overdrive_tone_s1_slavearbiterlockenable2 <= or_reduce(pio_overdrive_tone_s1_arb_share_counter_next_value);
  --cpu/data_master pio_overdrive_tone/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_overdrive_tone_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_overdrive_tone_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_overdrive_tone_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_overdrive_tone_s1 <= internal_cpu_data_master_requests_pio_overdrive_tone_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_overdrive_tone_s1_writedata mux, which is an e_mux
  pio_overdrive_tone_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_overdrive_tone_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_tone_s1;
  --cpu/data_master saved-grant pio_overdrive_tone/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_overdrive_tone_s1 <= internal_cpu_data_master_requests_pio_overdrive_tone_s1;
  --allow new arb cycle for pio_overdrive_tone/s1, which is an e_assign
  pio_overdrive_tone_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_overdrive_tone_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_overdrive_tone_s1_master_qreq_vector <= std_logic'('1');
  --pio_overdrive_tone_s1_reset_n assignment, which is an e_assign
  pio_overdrive_tone_s1_reset_n <= reset_n;
  pio_overdrive_tone_s1_chipselect <= internal_cpu_data_master_granted_pio_overdrive_tone_s1;
  --pio_overdrive_tone_s1_firsttransfer first transaction, which is an e_assign
  pio_overdrive_tone_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_overdrive_tone_s1_begins_xfer) = '1'), pio_overdrive_tone_s1_unreg_firsttransfer, pio_overdrive_tone_s1_reg_firsttransfer);
  --pio_overdrive_tone_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_overdrive_tone_s1_unreg_firsttransfer <= NOT ((pio_overdrive_tone_s1_slavearbiterlockenable AND pio_overdrive_tone_s1_any_continuerequest));
  --pio_overdrive_tone_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_tone_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_tone_s1_begins_xfer) = '1' then 
        pio_overdrive_tone_s1_reg_firsttransfer <= pio_overdrive_tone_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_overdrive_tone_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_overdrive_tone_s1_beginbursttransfer_internal <= pio_overdrive_tone_s1_begins_xfer;
  --~pio_overdrive_tone_s1_write_n assignment, which is an e_mux
  pio_overdrive_tone_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_overdrive_tone_s1 AND cpu_data_master_write));
  shifted_address_to_pio_overdrive_tone_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_overdrive_tone_s1_address mux, which is an e_mux
  pio_overdrive_tone_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_overdrive_tone_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_overdrive_tone_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_overdrive_tone_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_overdrive_tone_s1_end_xfer <= pio_overdrive_tone_s1_end_xfer;
    end if;

  end process;

  --pio_overdrive_tone_s1_waits_for_read in a cycle, which is an e_mux
  pio_overdrive_tone_s1_waits_for_read <= pio_overdrive_tone_s1_in_a_read_cycle AND pio_overdrive_tone_s1_begins_xfer;
  --pio_overdrive_tone_s1_in_a_read_cycle assignment, which is an e_assign
  pio_overdrive_tone_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_overdrive_tone_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_overdrive_tone_s1_in_a_read_cycle;
  --pio_overdrive_tone_s1_waits_for_write in a cycle, which is an e_mux
  pio_overdrive_tone_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_overdrive_tone_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_overdrive_tone_s1_in_a_write_cycle assignment, which is an e_assign
  pio_overdrive_tone_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_overdrive_tone_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_overdrive_tone_s1_in_a_write_cycle;
  wait_for_pio_overdrive_tone_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_overdrive_tone_s1 <= internal_cpu_data_master_granted_pio_overdrive_tone_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_overdrive_tone_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_tone_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_overdrive_tone_s1 <= internal_cpu_data_master_requests_pio_overdrive_tone_s1;
--synthesis translate_off
    --pio_overdrive_tone/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_overdrive_volume_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_overdrive_volume_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                 signal d1_pio_overdrive_volume_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_overdrive_volume_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_overdrive_volume_s1_chipselect : OUT STD_LOGIC;
                 signal pio_overdrive_volume_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_overdrive_volume_s1_reset_n : OUT STD_LOGIC;
                 signal pio_overdrive_volume_s1_write_n : OUT STD_LOGIC;
                 signal pio_overdrive_volume_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_overdrive_volume_s1_arbitrator;


architecture europa of pio_overdrive_volume_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal pio_overdrive_volume_s1_allgrants :  STD_LOGIC;
                signal pio_overdrive_volume_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_overdrive_volume_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_overdrive_volume_s1_any_continuerequest :  STD_LOGIC;
                signal pio_overdrive_volume_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_overdrive_volume_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_volume_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_volume_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_overdrive_volume_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_overdrive_volume_s1_begins_xfer :  STD_LOGIC;
                signal pio_overdrive_volume_s1_end_xfer :  STD_LOGIC;
                signal pio_overdrive_volume_s1_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_volume_s1_grant_vector :  STD_LOGIC;
                signal pio_overdrive_volume_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_overdrive_volume_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_overdrive_volume_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_overdrive_volume_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_overdrive_volume_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_volume_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_overdrive_volume_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_overdrive_volume_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_overdrive_volume_s1_waits_for_read :  STD_LOGIC;
                signal pio_overdrive_volume_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_overdrive_volume_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_overdrive_volume_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_overdrive_volume_s1_end_xfer;
    end if;

  end process;

  pio_overdrive_volume_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_overdrive_volume_s1);
  --assign pio_overdrive_volume_s1_readdata_from_sa = pio_overdrive_volume_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_overdrive_volume_s1_readdata_from_sa <= pio_overdrive_volume_s1_readdata;
  internal_cpu_data_master_requests_pio_overdrive_volume_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000000110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_overdrive_volume_s1_arb_share_counter set values, which is an e_mux
  pio_overdrive_volume_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_overdrive_volume_s1_non_bursting_master_requests mux, which is an e_mux
  pio_overdrive_volume_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_overdrive_volume_s1;
  --pio_overdrive_volume_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_overdrive_volume_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_overdrive_volume_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_overdrive_volume_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_overdrive_volume_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_volume_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_overdrive_volume_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_overdrive_volume_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_overdrive_volume_s1_allgrants all slave grants, which is an e_mux
  pio_overdrive_volume_s1_allgrants <= pio_overdrive_volume_s1_grant_vector;
  --pio_overdrive_volume_s1_end_xfer assignment, which is an e_assign
  pio_overdrive_volume_s1_end_xfer <= NOT ((pio_overdrive_volume_s1_waits_for_read OR pio_overdrive_volume_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_overdrive_volume_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_overdrive_volume_s1 <= pio_overdrive_volume_s1_end_xfer AND (((NOT pio_overdrive_volume_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_overdrive_volume_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_overdrive_volume_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_overdrive_volume_s1 AND pio_overdrive_volume_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_volume_s1 AND NOT pio_overdrive_volume_s1_non_bursting_master_requests));
  --pio_overdrive_volume_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_volume_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_volume_s1_arb_counter_enable) = '1' then 
        pio_overdrive_volume_s1_arb_share_counter <= pio_overdrive_volume_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_overdrive_volume_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_volume_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_overdrive_volume_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_overdrive_volume_s1)) OR ((end_xfer_arb_share_counter_term_pio_overdrive_volume_s1 AND NOT pio_overdrive_volume_s1_non_bursting_master_requests)))) = '1' then 
        pio_overdrive_volume_s1_slavearbiterlockenable <= or_reduce(pio_overdrive_volume_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_overdrive_volume/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_overdrive_volume_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_overdrive_volume_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_overdrive_volume_s1_slavearbiterlockenable2 <= or_reduce(pio_overdrive_volume_s1_arb_share_counter_next_value);
  --cpu/data_master pio_overdrive_volume/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_overdrive_volume_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_overdrive_volume_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_overdrive_volume_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_overdrive_volume_s1 <= internal_cpu_data_master_requests_pio_overdrive_volume_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_overdrive_volume_s1_writedata mux, which is an e_mux
  pio_overdrive_volume_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_overdrive_volume_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_volume_s1;
  --cpu/data_master saved-grant pio_overdrive_volume/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_overdrive_volume_s1 <= internal_cpu_data_master_requests_pio_overdrive_volume_s1;
  --allow new arb cycle for pio_overdrive_volume/s1, which is an e_assign
  pio_overdrive_volume_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_overdrive_volume_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_overdrive_volume_s1_master_qreq_vector <= std_logic'('1');
  --pio_overdrive_volume_s1_reset_n assignment, which is an e_assign
  pio_overdrive_volume_s1_reset_n <= reset_n;
  pio_overdrive_volume_s1_chipselect <= internal_cpu_data_master_granted_pio_overdrive_volume_s1;
  --pio_overdrive_volume_s1_firsttransfer first transaction, which is an e_assign
  pio_overdrive_volume_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_overdrive_volume_s1_begins_xfer) = '1'), pio_overdrive_volume_s1_unreg_firsttransfer, pio_overdrive_volume_s1_reg_firsttransfer);
  --pio_overdrive_volume_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_overdrive_volume_s1_unreg_firsttransfer <= NOT ((pio_overdrive_volume_s1_slavearbiterlockenable AND pio_overdrive_volume_s1_any_continuerequest));
  --pio_overdrive_volume_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_overdrive_volume_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_overdrive_volume_s1_begins_xfer) = '1' then 
        pio_overdrive_volume_s1_reg_firsttransfer <= pio_overdrive_volume_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_overdrive_volume_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_overdrive_volume_s1_beginbursttransfer_internal <= pio_overdrive_volume_s1_begins_xfer;
  --~pio_overdrive_volume_s1_write_n assignment, which is an e_mux
  pio_overdrive_volume_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_overdrive_volume_s1 AND cpu_data_master_write));
  shifted_address_to_pio_overdrive_volume_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_overdrive_volume_s1_address mux, which is an e_mux
  pio_overdrive_volume_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_overdrive_volume_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_overdrive_volume_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_overdrive_volume_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_overdrive_volume_s1_end_xfer <= pio_overdrive_volume_s1_end_xfer;
    end if;

  end process;

  --pio_overdrive_volume_s1_waits_for_read in a cycle, which is an e_mux
  pio_overdrive_volume_s1_waits_for_read <= pio_overdrive_volume_s1_in_a_read_cycle AND pio_overdrive_volume_s1_begins_xfer;
  --pio_overdrive_volume_s1_in_a_read_cycle assignment, which is an e_assign
  pio_overdrive_volume_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_overdrive_volume_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_overdrive_volume_s1_in_a_read_cycle;
  --pio_overdrive_volume_s1_waits_for_write in a cycle, which is an e_mux
  pio_overdrive_volume_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_overdrive_volume_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_overdrive_volume_s1_in_a_write_cycle assignment, which is an e_assign
  pio_overdrive_volume_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_overdrive_volume_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_overdrive_volume_s1_in_a_write_cycle;
  wait_for_pio_overdrive_volume_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_overdrive_volume_s1 <= internal_cpu_data_master_granted_pio_overdrive_volume_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_overdrive_volume_s1 <= internal_cpu_data_master_qualified_request_pio_overdrive_volume_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_overdrive_volume_s1 <= internal_cpu_data_master_requests_pio_overdrive_volume_s1;
--synthesis translate_off
    --pio_overdrive_volume/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_tremolo_stereo_bypass_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_tremolo_stereo_bypass_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                 signal d1_pio_tremolo_stereo_bypass_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_tremolo_stereo_bypass_s1_chipselect : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_bypass_s1_reset_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_bypass_s1_write_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_bypass_s1_writedata : OUT STD_LOGIC
              );
end entity pio_tremolo_stereo_bypass_s1_arbitrator;


architecture europa of pio_tremolo_stereo_bypass_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_allgrants :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_any_continuerequest :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_bypass_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_bypass_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_bypass_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_begins_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_end_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_grant_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_waits_for_read :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_tremolo_stereo_bypass_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_tremolo_stereo_bypass_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_tremolo_stereo_bypass_s1_end_xfer;
    end if;

  end process;

  pio_tremolo_stereo_bypass_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1);
  --assign pio_tremolo_stereo_bypass_s1_readdata_from_sa = pio_tremolo_stereo_bypass_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_tremolo_stereo_bypass_s1_readdata_from_sa <= pio_tremolo_stereo_bypass_s1_readdata;
  internal_cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000100110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_tremolo_stereo_bypass_s1_arb_share_counter set values, which is an e_mux
  pio_tremolo_stereo_bypass_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_tremolo_stereo_bypass_s1_non_bursting_master_requests mux, which is an e_mux
  pio_tremolo_stereo_bypass_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_tremolo_stereo_bypass_s1;
  --pio_tremolo_stereo_bypass_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_tremolo_stereo_bypass_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_tremolo_stereo_bypass_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_tremolo_stereo_bypass_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_tremolo_stereo_bypass_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_bypass_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_tremolo_stereo_bypass_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_bypass_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_tremolo_stereo_bypass_s1_allgrants all slave grants, which is an e_mux
  pio_tremolo_stereo_bypass_s1_allgrants <= pio_tremolo_stereo_bypass_s1_grant_vector;
  --pio_tremolo_stereo_bypass_s1_end_xfer assignment, which is an e_assign
  pio_tremolo_stereo_bypass_s1_end_xfer <= NOT ((pio_tremolo_stereo_bypass_s1_waits_for_read OR pio_tremolo_stereo_bypass_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_tremolo_stereo_bypass_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_tremolo_stereo_bypass_s1 <= pio_tremolo_stereo_bypass_s1_end_xfer AND (((NOT pio_tremolo_stereo_bypass_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_tremolo_stereo_bypass_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_tremolo_stereo_bypass_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_bypass_s1 AND pio_tremolo_stereo_bypass_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_bypass_s1 AND NOT pio_tremolo_stereo_bypass_s1_non_bursting_master_requests));
  --pio_tremolo_stereo_bypass_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_bypass_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_bypass_s1_arb_counter_enable) = '1' then 
        pio_tremolo_stereo_bypass_s1_arb_share_counter <= pio_tremolo_stereo_bypass_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_bypass_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_bypass_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_tremolo_stereo_bypass_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_tremolo_stereo_bypass_s1)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_bypass_s1 AND NOT pio_tremolo_stereo_bypass_s1_non_bursting_master_requests)))) = '1' then 
        pio_tremolo_stereo_bypass_s1_slavearbiterlockenable <= or_reduce(pio_tremolo_stereo_bypass_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_tremolo_stereo_bypass/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_tremolo_stereo_bypass_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_bypass_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_tremolo_stereo_bypass_s1_slavearbiterlockenable2 <= or_reduce(pio_tremolo_stereo_bypass_s1_arb_share_counter_next_value);
  --cpu/data_master pio_tremolo_stereo_bypass/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_tremolo_stereo_bypass_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_bypass_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_tremolo_stereo_bypass_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_tremolo_stereo_bypass_s1_writedata mux, which is an e_mux
  pio_tremolo_stereo_bypass_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1;
  --cpu/data_master saved-grant pio_tremolo_stereo_bypass/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_tremolo_stereo_bypass_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_bypass_s1;
  --allow new arb cycle for pio_tremolo_stereo_bypass/s1, which is an e_assign
  pio_tremolo_stereo_bypass_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_tremolo_stereo_bypass_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_tremolo_stereo_bypass_s1_master_qreq_vector <= std_logic'('1');
  --pio_tremolo_stereo_bypass_s1_reset_n assignment, which is an e_assign
  pio_tremolo_stereo_bypass_s1_reset_n <= reset_n;
  pio_tremolo_stereo_bypass_s1_chipselect <= internal_cpu_data_master_granted_pio_tremolo_stereo_bypass_s1;
  --pio_tremolo_stereo_bypass_s1_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_bypass_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_tremolo_stereo_bypass_s1_begins_xfer) = '1'), pio_tremolo_stereo_bypass_s1_unreg_firsttransfer, pio_tremolo_stereo_bypass_s1_reg_firsttransfer);
  --pio_tremolo_stereo_bypass_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_bypass_s1_unreg_firsttransfer <= NOT ((pio_tremolo_stereo_bypass_s1_slavearbiterlockenable AND pio_tremolo_stereo_bypass_s1_any_continuerequest));
  --pio_tremolo_stereo_bypass_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_bypass_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_bypass_s1_begins_xfer) = '1' then 
        pio_tremolo_stereo_bypass_s1_reg_firsttransfer <= pio_tremolo_stereo_bypass_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_bypass_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_tremolo_stereo_bypass_s1_beginbursttransfer_internal <= pio_tremolo_stereo_bypass_s1_begins_xfer;
  --~pio_tremolo_stereo_bypass_s1_write_n assignment, which is an e_mux
  pio_tremolo_stereo_bypass_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 AND cpu_data_master_write));
  shifted_address_to_pio_tremolo_stereo_bypass_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_tremolo_stereo_bypass_s1_address mux, which is an e_mux
  pio_tremolo_stereo_bypass_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_tremolo_stereo_bypass_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_tremolo_stereo_bypass_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_tremolo_stereo_bypass_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_tremolo_stereo_bypass_s1_end_xfer <= pio_tremolo_stereo_bypass_s1_end_xfer;
    end if;

  end process;

  --pio_tremolo_stereo_bypass_s1_waits_for_read in a cycle, which is an e_mux
  pio_tremolo_stereo_bypass_s1_waits_for_read <= pio_tremolo_stereo_bypass_s1_in_a_read_cycle AND pio_tremolo_stereo_bypass_s1_begins_xfer;
  --pio_tremolo_stereo_bypass_s1_in_a_read_cycle assignment, which is an e_assign
  pio_tremolo_stereo_bypass_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_tremolo_stereo_bypass_s1_in_a_read_cycle;
  --pio_tremolo_stereo_bypass_s1_waits_for_write in a cycle, which is an e_mux
  pio_tremolo_stereo_bypass_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_tremolo_stereo_bypass_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_tremolo_stereo_bypass_s1_in_a_write_cycle assignment, which is an e_assign
  pio_tremolo_stereo_bypass_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_tremolo_stereo_bypass_s1_in_a_write_cycle;
  wait_for_pio_tremolo_stereo_bypass_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 <= internal_cpu_data_master_granted_pio_tremolo_stereo_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_bypass_s1;
--synthesis translate_off
    --pio_tremolo_stereo_bypass/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_tremolo_stereo_depth_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_tremolo_stereo_depth_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                 signal d1_pio_tremolo_stereo_depth_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_depth_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_tremolo_stereo_depth_s1_chipselect : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_depth_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pio_tremolo_stereo_depth_s1_reset_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_depth_s1_write_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_depth_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pio_tremolo_stereo_depth_s1_arbitrator;


architecture europa of pio_tremolo_stereo_depth_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_allgrants :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_any_continuerequest :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_depth_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_depth_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_depth_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_begins_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_end_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_grant_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_waits_for_read :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_tremolo_stereo_depth_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_tremolo_stereo_depth_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_tremolo_stereo_depth_s1_end_xfer;
    end if;

  end process;

  pio_tremolo_stereo_depth_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1);
  --assign pio_tremolo_stereo_depth_s1_readdata_from_sa = pio_tremolo_stereo_depth_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_tremolo_stereo_depth_s1_readdata_from_sa <= pio_tremolo_stereo_depth_s1_readdata;
  internal_cpu_data_master_requests_pio_tremolo_stereo_depth_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000101000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_tremolo_stereo_depth_s1_arb_share_counter set values, which is an e_mux
  pio_tremolo_stereo_depth_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_tremolo_stereo_depth_s1_non_bursting_master_requests mux, which is an e_mux
  pio_tremolo_stereo_depth_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_tremolo_stereo_depth_s1;
  --pio_tremolo_stereo_depth_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_tremolo_stereo_depth_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_tremolo_stereo_depth_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_tremolo_stereo_depth_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_tremolo_stereo_depth_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_depth_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_tremolo_stereo_depth_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_depth_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_tremolo_stereo_depth_s1_allgrants all slave grants, which is an e_mux
  pio_tremolo_stereo_depth_s1_allgrants <= pio_tremolo_stereo_depth_s1_grant_vector;
  --pio_tremolo_stereo_depth_s1_end_xfer assignment, which is an e_assign
  pio_tremolo_stereo_depth_s1_end_xfer <= NOT ((pio_tremolo_stereo_depth_s1_waits_for_read OR pio_tremolo_stereo_depth_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_tremolo_stereo_depth_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_tremolo_stereo_depth_s1 <= pio_tremolo_stereo_depth_s1_end_xfer AND (((NOT pio_tremolo_stereo_depth_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_tremolo_stereo_depth_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_tremolo_stereo_depth_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_depth_s1 AND pio_tremolo_stereo_depth_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_depth_s1 AND NOT pio_tremolo_stereo_depth_s1_non_bursting_master_requests));
  --pio_tremolo_stereo_depth_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_depth_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_depth_s1_arb_counter_enable) = '1' then 
        pio_tremolo_stereo_depth_s1_arb_share_counter <= pio_tremolo_stereo_depth_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_depth_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_depth_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_tremolo_stereo_depth_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_tremolo_stereo_depth_s1)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_depth_s1 AND NOT pio_tremolo_stereo_depth_s1_non_bursting_master_requests)))) = '1' then 
        pio_tremolo_stereo_depth_s1_slavearbiterlockenable <= or_reduce(pio_tremolo_stereo_depth_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_tremolo_stereo_depth/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_tremolo_stereo_depth_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_depth_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_tremolo_stereo_depth_s1_slavearbiterlockenable2 <= or_reduce(pio_tremolo_stereo_depth_s1_arb_share_counter_next_value);
  --cpu/data_master pio_tremolo_stereo_depth/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_tremolo_stereo_depth_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_depth_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_tremolo_stereo_depth_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_depth_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_tremolo_stereo_depth_s1_writedata mux, which is an e_mux
  pio_tremolo_stereo_depth_s1_writedata <= cpu_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_tremolo_stereo_depth_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1;
  --cpu/data_master saved-grant pio_tremolo_stereo_depth/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_tremolo_stereo_depth_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_depth_s1;
  --allow new arb cycle for pio_tremolo_stereo_depth/s1, which is an e_assign
  pio_tremolo_stereo_depth_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_tremolo_stereo_depth_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_tremolo_stereo_depth_s1_master_qreq_vector <= std_logic'('1');
  --pio_tremolo_stereo_depth_s1_reset_n assignment, which is an e_assign
  pio_tremolo_stereo_depth_s1_reset_n <= reset_n;
  pio_tremolo_stereo_depth_s1_chipselect <= internal_cpu_data_master_granted_pio_tremolo_stereo_depth_s1;
  --pio_tremolo_stereo_depth_s1_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_depth_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_tremolo_stereo_depth_s1_begins_xfer) = '1'), pio_tremolo_stereo_depth_s1_unreg_firsttransfer, pio_tremolo_stereo_depth_s1_reg_firsttransfer);
  --pio_tremolo_stereo_depth_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_depth_s1_unreg_firsttransfer <= NOT ((pio_tremolo_stereo_depth_s1_slavearbiterlockenable AND pio_tremolo_stereo_depth_s1_any_continuerequest));
  --pio_tremolo_stereo_depth_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_depth_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_depth_s1_begins_xfer) = '1' then 
        pio_tremolo_stereo_depth_s1_reg_firsttransfer <= pio_tremolo_stereo_depth_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_depth_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_tremolo_stereo_depth_s1_beginbursttransfer_internal <= pio_tremolo_stereo_depth_s1_begins_xfer;
  --~pio_tremolo_stereo_depth_s1_write_n assignment, which is an e_mux
  pio_tremolo_stereo_depth_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_tremolo_stereo_depth_s1 AND cpu_data_master_write));
  shifted_address_to_pio_tremolo_stereo_depth_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_tremolo_stereo_depth_s1_address mux, which is an e_mux
  pio_tremolo_stereo_depth_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_tremolo_stereo_depth_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_tremolo_stereo_depth_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_tremolo_stereo_depth_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_tremolo_stereo_depth_s1_end_xfer <= pio_tremolo_stereo_depth_s1_end_xfer;
    end if;

  end process;

  --pio_tremolo_stereo_depth_s1_waits_for_read in a cycle, which is an e_mux
  pio_tremolo_stereo_depth_s1_waits_for_read <= pio_tremolo_stereo_depth_s1_in_a_read_cycle AND pio_tremolo_stereo_depth_s1_begins_xfer;
  --pio_tremolo_stereo_depth_s1_in_a_read_cycle assignment, which is an e_assign
  pio_tremolo_stereo_depth_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_depth_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_tremolo_stereo_depth_s1_in_a_read_cycle;
  --pio_tremolo_stereo_depth_s1_waits_for_write in a cycle, which is an e_mux
  pio_tremolo_stereo_depth_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_tremolo_stereo_depth_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_tremolo_stereo_depth_s1_in_a_write_cycle assignment, which is an e_assign
  pio_tremolo_stereo_depth_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_depth_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_tremolo_stereo_depth_s1_in_a_write_cycle;
  wait_for_pio_tremolo_stereo_depth_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_tremolo_stereo_depth_s1 <= internal_cpu_data_master_granted_pio_tremolo_stereo_depth_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_tremolo_stereo_depth_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_depth_s1;
--synthesis translate_off
    --pio_tremolo_stereo_depth/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_tremolo_stereo_mode_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_tremolo_stereo_mode_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                 signal d1_pio_tremolo_stereo_mode_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_mode_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_tremolo_stereo_mode_s1_chipselect : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_mode_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_mode_s1_reset_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_mode_s1_write_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_mode_s1_writedata : OUT STD_LOGIC
              );
end entity pio_tremolo_stereo_mode_s1_arbitrator;


architecture europa of pio_tremolo_stereo_mode_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_allgrants :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_any_continuerequest :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_mode_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_mode_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_mode_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_begins_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_end_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_grant_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_waits_for_read :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_tremolo_stereo_mode_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_tremolo_stereo_mode_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_tremolo_stereo_mode_s1_end_xfer;
    end if;

  end process;

  pio_tremolo_stereo_mode_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1);
  --assign pio_tremolo_stereo_mode_s1_readdata_from_sa = pio_tremolo_stereo_mode_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_tremolo_stereo_mode_s1_readdata_from_sa <= pio_tremolo_stereo_mode_s1_readdata;
  internal_cpu_data_master_requests_pio_tremolo_stereo_mode_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110000000000000000010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_tremolo_stereo_mode_s1_arb_share_counter set values, which is an e_mux
  pio_tremolo_stereo_mode_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_tremolo_stereo_mode_s1_non_bursting_master_requests mux, which is an e_mux
  pio_tremolo_stereo_mode_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_tremolo_stereo_mode_s1;
  --pio_tremolo_stereo_mode_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_tremolo_stereo_mode_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_tremolo_stereo_mode_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_tremolo_stereo_mode_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_tremolo_stereo_mode_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_mode_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_tremolo_stereo_mode_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_mode_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_tremolo_stereo_mode_s1_allgrants all slave grants, which is an e_mux
  pio_tremolo_stereo_mode_s1_allgrants <= pio_tremolo_stereo_mode_s1_grant_vector;
  --pio_tremolo_stereo_mode_s1_end_xfer assignment, which is an e_assign
  pio_tremolo_stereo_mode_s1_end_xfer <= NOT ((pio_tremolo_stereo_mode_s1_waits_for_read OR pio_tremolo_stereo_mode_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_tremolo_stereo_mode_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_tremolo_stereo_mode_s1 <= pio_tremolo_stereo_mode_s1_end_xfer AND (((NOT pio_tremolo_stereo_mode_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_tremolo_stereo_mode_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_tremolo_stereo_mode_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_mode_s1 AND pio_tremolo_stereo_mode_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_mode_s1 AND NOT pio_tremolo_stereo_mode_s1_non_bursting_master_requests));
  --pio_tremolo_stereo_mode_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_mode_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_mode_s1_arb_counter_enable) = '1' then 
        pio_tremolo_stereo_mode_s1_arb_share_counter <= pio_tremolo_stereo_mode_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_mode_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_mode_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_tremolo_stereo_mode_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_tremolo_stereo_mode_s1)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_mode_s1 AND NOT pio_tremolo_stereo_mode_s1_non_bursting_master_requests)))) = '1' then 
        pio_tremolo_stereo_mode_s1_slavearbiterlockenable <= or_reduce(pio_tremolo_stereo_mode_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_tremolo_stereo_mode/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_tremolo_stereo_mode_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_mode_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_tremolo_stereo_mode_s1_slavearbiterlockenable2 <= or_reduce(pio_tremolo_stereo_mode_s1_arb_share_counter_next_value);
  --cpu/data_master pio_tremolo_stereo_mode/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_tremolo_stereo_mode_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_mode_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_tremolo_stereo_mode_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_mode_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_tremolo_stereo_mode_s1_writedata mux, which is an e_mux
  pio_tremolo_stereo_mode_s1_writedata <= cpu_data_master_writedata(0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_tremolo_stereo_mode_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1;
  --cpu/data_master saved-grant pio_tremolo_stereo_mode/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_tremolo_stereo_mode_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_mode_s1;
  --allow new arb cycle for pio_tremolo_stereo_mode/s1, which is an e_assign
  pio_tremolo_stereo_mode_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_tremolo_stereo_mode_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_tremolo_stereo_mode_s1_master_qreq_vector <= std_logic'('1');
  --pio_tremolo_stereo_mode_s1_reset_n assignment, which is an e_assign
  pio_tremolo_stereo_mode_s1_reset_n <= reset_n;
  pio_tremolo_stereo_mode_s1_chipselect <= internal_cpu_data_master_granted_pio_tremolo_stereo_mode_s1;
  --pio_tremolo_stereo_mode_s1_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_mode_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_tremolo_stereo_mode_s1_begins_xfer) = '1'), pio_tremolo_stereo_mode_s1_unreg_firsttransfer, pio_tremolo_stereo_mode_s1_reg_firsttransfer);
  --pio_tremolo_stereo_mode_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_mode_s1_unreg_firsttransfer <= NOT ((pio_tremolo_stereo_mode_s1_slavearbiterlockenable AND pio_tremolo_stereo_mode_s1_any_continuerequest));
  --pio_tremolo_stereo_mode_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_mode_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_mode_s1_begins_xfer) = '1' then 
        pio_tremolo_stereo_mode_s1_reg_firsttransfer <= pio_tremolo_stereo_mode_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_mode_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_tremolo_stereo_mode_s1_beginbursttransfer_internal <= pio_tremolo_stereo_mode_s1_begins_xfer;
  --~pio_tremolo_stereo_mode_s1_write_n assignment, which is an e_mux
  pio_tremolo_stereo_mode_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_tremolo_stereo_mode_s1 AND cpu_data_master_write));
  shifted_address_to_pio_tremolo_stereo_mode_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_tremolo_stereo_mode_s1_address mux, which is an e_mux
  pio_tremolo_stereo_mode_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_tremolo_stereo_mode_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_tremolo_stereo_mode_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_tremolo_stereo_mode_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_tremolo_stereo_mode_s1_end_xfer <= pio_tremolo_stereo_mode_s1_end_xfer;
    end if;

  end process;

  --pio_tremolo_stereo_mode_s1_waits_for_read in a cycle, which is an e_mux
  pio_tremolo_stereo_mode_s1_waits_for_read <= pio_tremolo_stereo_mode_s1_in_a_read_cycle AND pio_tremolo_stereo_mode_s1_begins_xfer;
  --pio_tremolo_stereo_mode_s1_in_a_read_cycle assignment, which is an e_assign
  pio_tremolo_stereo_mode_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_mode_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_tremolo_stereo_mode_s1_in_a_read_cycle;
  --pio_tremolo_stereo_mode_s1_waits_for_write in a cycle, which is an e_mux
  pio_tremolo_stereo_mode_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_tremolo_stereo_mode_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_tremolo_stereo_mode_s1_in_a_write_cycle assignment, which is an e_assign
  pio_tremolo_stereo_mode_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_mode_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_tremolo_stereo_mode_s1_in_a_write_cycle;
  wait_for_pio_tremolo_stereo_mode_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_tremolo_stereo_mode_s1 <= internal_cpu_data_master_granted_pio_tremolo_stereo_mode_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_tremolo_stereo_mode_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_mode_s1;
--synthesis translate_off
    --pio_tremolo_stereo_mode/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_tremolo_stereo_sweep_a_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_tremolo_stereo_sweep_a_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                 signal d1_pio_tremolo_stereo_sweep_a_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_a_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_tremolo_stereo_sweep_a_s1_chipselect : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_a_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pio_tremolo_stereo_sweep_a_s1_reset_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_a_s1_write_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_a_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
              );
end entity pio_tremolo_stereo_sweep_a_s1_arbitrator;


architecture europa of pio_tremolo_stereo_sweep_a_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_allgrants :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_any_continuerequest :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_a_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_a_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_a_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_begins_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_end_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_grant_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_waits_for_read :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_tremolo_stereo_sweep_a_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_tremolo_stereo_sweep_a_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_tremolo_stereo_sweep_a_s1_end_xfer;
    end if;

  end process;

  pio_tremolo_stereo_sweep_a_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1);
  --assign pio_tremolo_stereo_sweep_a_s1_readdata_from_sa = pio_tremolo_stereo_sweep_a_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_readdata_from_sa <= pio_tremolo_stereo_sweep_a_s1_readdata;
  internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000101010000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_tremolo_stereo_sweep_a_s1_arb_share_counter set values, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_tremolo_stereo_sweep_a_s1_non_bursting_master_requests mux, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1;
  --pio_tremolo_stereo_sweep_a_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_tremolo_stereo_sweep_a_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_tremolo_stereo_sweep_a_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_sweep_a_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_tremolo_stereo_sweep_a_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_sweep_a_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_tremolo_stereo_sweep_a_s1_allgrants all slave grants, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_allgrants <= pio_tremolo_stereo_sweep_a_s1_grant_vector;
  --pio_tremolo_stereo_sweep_a_s1_end_xfer assignment, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_end_xfer <= NOT ((pio_tremolo_stereo_sweep_a_s1_waits_for_read OR pio_tremolo_stereo_sweep_a_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_a_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_a_s1 <= pio_tremolo_stereo_sweep_a_s1_end_xfer AND (((NOT pio_tremolo_stereo_sweep_a_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_tremolo_stereo_sweep_a_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_a_s1 AND pio_tremolo_stereo_sweep_a_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_a_s1 AND NOT pio_tremolo_stereo_sweep_a_s1_non_bursting_master_requests));
  --pio_tremolo_stereo_sweep_a_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_sweep_a_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_sweep_a_s1_arb_counter_enable) = '1' then 
        pio_tremolo_stereo_sweep_a_s1_arb_share_counter <= pio_tremolo_stereo_sweep_a_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_tremolo_stereo_sweep_a_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_a_s1)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_a_s1 AND NOT pio_tremolo_stereo_sweep_a_s1_non_bursting_master_requests)))) = '1' then 
        pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable <= or_reduce(pio_tremolo_stereo_sweep_a_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_tremolo_stereo_sweep_a/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable2 <= or_reduce(pio_tremolo_stereo_sweep_a_s1_arb_share_counter_next_value);
  --cpu/data_master pio_tremolo_stereo_sweep_a/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_sweep_a_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_tremolo_stereo_sweep_a_s1_writedata mux, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_writedata <= cpu_data_master_writedata (3 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1;
  --cpu/data_master saved-grant pio_tremolo_stereo_sweep_a/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_tremolo_stereo_sweep_a_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1;
  --allow new arb cycle for pio_tremolo_stereo_sweep_a/s1, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_tremolo_stereo_sweep_a_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_tremolo_stereo_sweep_a_s1_master_qreq_vector <= std_logic'('1');
  --pio_tremolo_stereo_sweep_a_s1_reset_n assignment, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_reset_n <= reset_n;
  pio_tremolo_stereo_sweep_a_s1_chipselect <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1;
  --pio_tremolo_stereo_sweep_a_s1_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_tremolo_stereo_sweep_a_s1_begins_xfer) = '1'), pio_tremolo_stereo_sweep_a_s1_unreg_firsttransfer, pio_tremolo_stereo_sweep_a_s1_reg_firsttransfer);
  --pio_tremolo_stereo_sweep_a_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_unreg_firsttransfer <= NOT ((pio_tremolo_stereo_sweep_a_s1_slavearbiterlockenable AND pio_tremolo_stereo_sweep_a_s1_any_continuerequest));
  --pio_tremolo_stereo_sweep_a_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_sweep_a_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_sweep_a_s1_begins_xfer) = '1' then 
        pio_tremolo_stereo_sweep_a_s1_reg_firsttransfer <= pio_tremolo_stereo_sweep_a_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_sweep_a_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_beginbursttransfer_internal <= pio_tremolo_stereo_sweep_a_s1_begins_xfer;
  --~pio_tremolo_stereo_sweep_a_s1_write_n assignment, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 AND cpu_data_master_write));
  shifted_address_to_pio_tremolo_stereo_sweep_a_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_tremolo_stereo_sweep_a_s1_address mux, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_tremolo_stereo_sweep_a_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_tremolo_stereo_sweep_a_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_tremolo_stereo_sweep_a_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_tremolo_stereo_sweep_a_s1_end_xfer <= pio_tremolo_stereo_sweep_a_s1_end_xfer;
    end if;

  end process;

  --pio_tremolo_stereo_sweep_a_s1_waits_for_read in a cycle, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_waits_for_read <= pio_tremolo_stereo_sweep_a_s1_in_a_read_cycle AND pio_tremolo_stereo_sweep_a_s1_begins_xfer;
  --pio_tremolo_stereo_sweep_a_s1_in_a_read_cycle assignment, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_tremolo_stereo_sweep_a_s1_in_a_read_cycle;
  --pio_tremolo_stereo_sweep_a_s1_waits_for_write in a cycle, which is an e_mux
  pio_tremolo_stereo_sweep_a_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_tremolo_stereo_sweep_a_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_tremolo_stereo_sweep_a_s1_in_a_write_cycle assignment, which is an e_assign
  pio_tremolo_stereo_sweep_a_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_tremolo_stereo_sweep_a_s1_in_a_write_cycle;
  wait_for_pio_tremolo_stereo_sweep_a_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1;
--synthesis translate_off
    --pio_tremolo_stereo_sweep_a/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pio_tremolo_stereo_sweep_b_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pio_tremolo_stereo_sweep_b_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                 signal d1_pio_tremolo_stereo_sweep_b_s1_end_xfer : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_b_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pio_tremolo_stereo_sweep_b_s1_chipselect : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_b_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pio_tremolo_stereo_sweep_b_s1_reset_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_b_s1_write_n : OUT STD_LOGIC;
                 signal pio_tremolo_stereo_sweep_b_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
              );
end entity pio_tremolo_stereo_sweep_b_s1_arbitrator;


architecture europa of pio_tremolo_stereo_sweep_b_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_allgrants :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_any_continuerequest :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_arb_counter_enable :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_b_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_b_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_b_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_begins_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_end_xfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_grant_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_in_a_read_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_in_a_write_cycle :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_master_qreq_vector :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_reg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_waits_for_read :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pio_tremolo_stereo_sweep_b_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pio_tremolo_stereo_sweep_b_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pio_tremolo_stereo_sweep_b_s1_end_xfer;
    end if;

  end process;

  pio_tremolo_stereo_sweep_b_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1);
  --assign pio_tremolo_stereo_sweep_b_s1_readdata_from_sa = pio_tremolo_stereo_sweep_b_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_readdata_from_sa <= pio_tremolo_stereo_sweep_b_s1_readdata;
  internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --pio_tremolo_stereo_sweep_b_s1_arb_share_counter set values, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_arb_share_set_values <= std_logic_vector'("001");
  --pio_tremolo_stereo_sweep_b_s1_non_bursting_master_requests mux, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1;
  --pio_tremolo_stereo_sweep_b_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pio_tremolo_stereo_sweep_b_s1_arb_share_counter_next_value assignment, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pio_tremolo_stereo_sweep_b_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_sweep_b_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pio_tremolo_stereo_sweep_b_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pio_tremolo_stereo_sweep_b_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pio_tremolo_stereo_sweep_b_s1_allgrants all slave grants, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_allgrants <= pio_tremolo_stereo_sweep_b_s1_grant_vector;
  --pio_tremolo_stereo_sweep_b_s1_end_xfer assignment, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_end_xfer <= NOT ((pio_tremolo_stereo_sweep_b_s1_waits_for_read OR pio_tremolo_stereo_sweep_b_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_b_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_b_s1 <= pio_tremolo_stereo_sweep_b_s1_end_xfer AND (((NOT pio_tremolo_stereo_sweep_b_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pio_tremolo_stereo_sweep_b_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_b_s1 AND pio_tremolo_stereo_sweep_b_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_b_s1 AND NOT pio_tremolo_stereo_sweep_b_s1_non_bursting_master_requests));
  --pio_tremolo_stereo_sweep_b_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_sweep_b_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_sweep_b_s1_arb_counter_enable) = '1' then 
        pio_tremolo_stereo_sweep_b_s1_arb_share_counter <= pio_tremolo_stereo_sweep_b_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pio_tremolo_stereo_sweep_b_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_b_s1)) OR ((end_xfer_arb_share_counter_term_pio_tremolo_stereo_sweep_b_s1 AND NOT pio_tremolo_stereo_sweep_b_s1_non_bursting_master_requests)))) = '1' then 
        pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable <= or_reduce(pio_tremolo_stereo_sweep_b_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pio_tremolo_stereo_sweep_b/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable2 <= or_reduce(pio_tremolo_stereo_sweep_b_s1_arb_share_counter_next_value);
  --cpu/data_master pio_tremolo_stereo_sweep_b/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pio_tremolo_stereo_sweep_b_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 AND NOT (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write));
  --pio_tremolo_stereo_sweep_b_s1_writedata mux, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_writedata <= cpu_data_master_writedata (3 DOWNTO 0);
  --master is always granted when requested
  internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1;
  --cpu/data_master saved-grant pio_tremolo_stereo_sweep_b/s1, which is an e_assign
  cpu_data_master_saved_grant_pio_tremolo_stereo_sweep_b_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1;
  --allow new arb cycle for pio_tremolo_stereo_sweep_b/s1, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pio_tremolo_stereo_sweep_b_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pio_tremolo_stereo_sweep_b_s1_master_qreq_vector <= std_logic'('1');
  --pio_tremolo_stereo_sweep_b_s1_reset_n assignment, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_reset_n <= reset_n;
  pio_tremolo_stereo_sweep_b_s1_chipselect <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1;
  --pio_tremolo_stereo_sweep_b_s1_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pio_tremolo_stereo_sweep_b_s1_begins_xfer) = '1'), pio_tremolo_stereo_sweep_b_s1_unreg_firsttransfer, pio_tremolo_stereo_sweep_b_s1_reg_firsttransfer);
  --pio_tremolo_stereo_sweep_b_s1_unreg_firsttransfer first transaction, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_unreg_firsttransfer <= NOT ((pio_tremolo_stereo_sweep_b_s1_slavearbiterlockenable AND pio_tremolo_stereo_sweep_b_s1_any_continuerequest));
  --pio_tremolo_stereo_sweep_b_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pio_tremolo_stereo_sweep_b_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pio_tremolo_stereo_sweep_b_s1_begins_xfer) = '1' then 
        pio_tremolo_stereo_sweep_b_s1_reg_firsttransfer <= pio_tremolo_stereo_sweep_b_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pio_tremolo_stereo_sweep_b_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_beginbursttransfer_internal <= pio_tremolo_stereo_sweep_b_s1_begins_xfer;
  --~pio_tremolo_stereo_sweep_b_s1_write_n assignment, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_write_n <= NOT ((internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 AND cpu_data_master_write));
  shifted_address_to_pio_tremolo_stereo_sweep_b_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pio_tremolo_stereo_sweep_b_s1_address mux, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_address <= A_EXT (A_SRL(shifted_address_to_pio_tremolo_stereo_sweep_b_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pio_tremolo_stereo_sweep_b_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pio_tremolo_stereo_sweep_b_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pio_tremolo_stereo_sweep_b_s1_end_xfer <= pio_tremolo_stereo_sweep_b_s1_end_xfer;
    end if;

  end process;

  --pio_tremolo_stereo_sweep_b_s1_waits_for_read in a cycle, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_waits_for_read <= pio_tremolo_stereo_sweep_b_s1_in_a_read_cycle AND pio_tremolo_stereo_sweep_b_s1_begins_xfer;
  --pio_tremolo_stereo_sweep_b_s1_in_a_read_cycle assignment, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_in_a_read_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pio_tremolo_stereo_sweep_b_s1_in_a_read_cycle;
  --pio_tremolo_stereo_sweep_b_s1_waits_for_write in a cycle, which is an e_mux
  pio_tremolo_stereo_sweep_b_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pio_tremolo_stereo_sweep_b_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pio_tremolo_stereo_sweep_b_s1_in_a_write_cycle assignment, which is an e_assign
  pio_tremolo_stereo_sweep_b_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pio_tremolo_stereo_sweep_b_s1_in_a_write_cycle;
  wait_for_pio_tremolo_stereo_sweep_b_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 <= internal_cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 <= internal_cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 <= internal_cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1;
--synthesis translate_off
    --pio_tremolo_stereo_sweep_b/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pixel_buffer_avalon_pixel_buffer_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                 signal d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_slave_read : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_slave_reset : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_slave_write : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC
              );
end entity pixel_buffer_avalon_pixel_buffer_slave_arbitrator;


architecture europa of pixel_buffer_avalon_pixel_buffer_slave_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_allgrants :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_any_continuerequest :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_arb_counter_enable :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_begins_xfer :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_end_xfer :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_firsttransfer :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_grant_vector :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_in_a_read_cycle :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_in_a_write_cycle :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_master_qreq_vector :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_non_bursting_master_requests :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_reg_firsttransfer :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_unreg_firsttransfer :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_waits_for_read :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pixel_buffer_avalon_pixel_buffer_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_pixel_buffer_avalon_pixel_buffer_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pixel_buffer_avalon_pixel_buffer_slave_end_xfer;
    end if;

  end process;

  pixel_buffer_avalon_pixel_buffer_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave);
  --assign pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa = pixel_buffer_avalon_pixel_buffer_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa <= pixel_buffer_avalon_pixel_buffer_slave_readdata;
  internal_cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("110100000011000000100000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --registered rdv signal_name registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave assignment, which is an e_assign
  registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave <= cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register_in;
  --pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter set values, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_arb_share_set_values <= std_logic_vector'("001");
  --pixel_buffer_avalon_pixel_buffer_slave_non_bursting_master_requests mux, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave;
  --pixel_buffer_avalon_pixel_buffer_slave_any_bursting_master_saved_grant mux, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter_next_value assignment, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pixel_buffer_avalon_pixel_buffer_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pixel_buffer_avalon_pixel_buffer_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --pixel_buffer_avalon_pixel_buffer_slave_allgrants all slave grants, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_allgrants <= pixel_buffer_avalon_pixel_buffer_slave_grant_vector;
  --pixel_buffer_avalon_pixel_buffer_slave_end_xfer assignment, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_end_xfer <= NOT ((pixel_buffer_avalon_pixel_buffer_slave_waits_for_read OR pixel_buffer_avalon_pixel_buffer_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_pixel_buffer_avalon_pixel_buffer_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pixel_buffer_avalon_pixel_buffer_slave <= pixel_buffer_avalon_pixel_buffer_slave_end_xfer AND (((NOT pixel_buffer_avalon_pixel_buffer_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter arbitration counter enable, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pixel_buffer_avalon_pixel_buffer_slave AND pixel_buffer_avalon_pixel_buffer_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_pixel_buffer_avalon_pixel_buffer_slave AND NOT pixel_buffer_avalon_pixel_buffer_slave_non_bursting_master_requests));
  --pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(pixel_buffer_avalon_pixel_buffer_slave_arb_counter_enable) = '1' then 
        pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter <= pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pixel_buffer_avalon_pixel_buffer_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_pixel_buffer_avalon_pixel_buffer_slave)) OR ((end_xfer_arb_share_counter_term_pixel_buffer_avalon_pixel_buffer_slave AND NOT pixel_buffer_avalon_pixel_buffer_slave_non_bursting_master_requests)))) = '1' then 
        pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable <= or_reduce(pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master pixel_buffer/avalon_pixel_buffer_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable2 <= or_reduce(pixel_buffer_avalon_pixel_buffer_slave_arb_share_counter_next_value);
  --cpu/data_master pixel_buffer/avalon_pixel_buffer_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --pixel_buffer_avalon_pixel_buffer_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave <= internal_cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave AND NOT ((((cpu_data_master_read AND (cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register))) OR (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write))));
  --cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register_in <= ((internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave AND cpu_data_master_read) AND NOT pixel_buffer_avalon_pixel_buffer_slave_waits_for_read) AND NOT (cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register);
  --shift register p1 cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register) & A_ToStdLogicVector(cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register_in)));
  --cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register <= p1_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave, which is an e_mux
  cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave <= cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave_shift_register;
  --pixel_buffer_avalon_pixel_buffer_slave_writedata mux, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave <= internal_cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave;
  --cpu/data_master saved-grant pixel_buffer/avalon_pixel_buffer_slave, which is an e_assign
  cpu_data_master_saved_grant_pixel_buffer_avalon_pixel_buffer_slave <= internal_cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave;
  --allow new arb cycle for pixel_buffer/avalon_pixel_buffer_slave, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pixel_buffer_avalon_pixel_buffer_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pixel_buffer_avalon_pixel_buffer_slave_master_qreq_vector <= std_logic'('1');
  --~pixel_buffer_avalon_pixel_buffer_slave_reset assignment, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_reset <= NOT reset_n;
  --pixel_buffer_avalon_pixel_buffer_slave_firsttransfer first transaction, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_firsttransfer <= A_WE_StdLogic((std_logic'(pixel_buffer_avalon_pixel_buffer_slave_begins_xfer) = '1'), pixel_buffer_avalon_pixel_buffer_slave_unreg_firsttransfer, pixel_buffer_avalon_pixel_buffer_slave_reg_firsttransfer);
  --pixel_buffer_avalon_pixel_buffer_slave_unreg_firsttransfer first transaction, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_unreg_firsttransfer <= NOT ((pixel_buffer_avalon_pixel_buffer_slave_slavearbiterlockenable AND pixel_buffer_avalon_pixel_buffer_slave_any_continuerequest));
  --pixel_buffer_avalon_pixel_buffer_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pixel_buffer_avalon_pixel_buffer_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pixel_buffer_avalon_pixel_buffer_slave_begins_xfer) = '1' then 
        pixel_buffer_avalon_pixel_buffer_slave_reg_firsttransfer <= pixel_buffer_avalon_pixel_buffer_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pixel_buffer_avalon_pixel_buffer_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_beginbursttransfer_internal <= pixel_buffer_avalon_pixel_buffer_slave_begins_xfer;
  --pixel_buffer_avalon_pixel_buffer_slave_read assignment, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_read <= internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave AND cpu_data_master_read;
  --pixel_buffer_avalon_pixel_buffer_slave_write assignment, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_write <= internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave AND cpu_data_master_write;
  shifted_address_to_pixel_buffer_avalon_pixel_buffer_slave_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pixel_buffer_avalon_pixel_buffer_slave_address mux, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_address <= A_EXT (A_SRL(shifted_address_to_pixel_buffer_avalon_pixel_buffer_slave_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer <= pixel_buffer_avalon_pixel_buffer_slave_end_xfer;
    end if;

  end process;

  --pixel_buffer_avalon_pixel_buffer_slave_waits_for_read in a cycle, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pixel_buffer_avalon_pixel_buffer_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pixel_buffer_avalon_pixel_buffer_slave_in_a_read_cycle assignment, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_in_a_read_cycle <= internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pixel_buffer_avalon_pixel_buffer_slave_in_a_read_cycle;
  --pixel_buffer_avalon_pixel_buffer_slave_waits_for_write in a cycle, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pixel_buffer_avalon_pixel_buffer_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pixel_buffer_avalon_pixel_buffer_slave_in_a_write_cycle assignment, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_slave_in_a_write_cycle <= internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pixel_buffer_avalon_pixel_buffer_slave_in_a_write_cycle;
  wait_for_pixel_buffer_avalon_pixel_buffer_slave_counter <= std_logic'('0');
  --pixel_buffer_avalon_pixel_buffer_slave_byteenable byte enable port mux, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave <= internal_cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave <= internal_cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave <= internal_cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave;
--synthesis translate_off
    --pixel_buffer/avalon_pixel_buffer_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pixel_buffer_avalon_pixel_buffer_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_read : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal pixel_buffer_avalon_pixel_buffer_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_master_latency_counter : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_master_readdatavalid : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_waitrequest : OUT STD_LOGIC
              );
end entity pixel_buffer_avalon_pixel_buffer_master_arbitrator;


architecture europa of pixel_buffer_avalon_pixel_buffer_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_pixel_buffer_avalon_pixel_buffer_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_pixel_buffer_avalon_pixel_buffer_master_latency_counter :  STD_LOGIC;
                signal internal_pixel_buffer_avalon_pixel_buffer_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_pixel_buffer_avalon_pixel_buffer_master_latency_counter :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_master_is_granted_some_slave :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_read_but_no_slave_selected :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_read_last_time :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_run :  STD_LOGIC;
                signal pre_flush_pixel_buffer_avalon_pixel_buffer_master_readdatavalid :  STD_LOGIC;
                signal r_7 :  STD_LOGIC;

begin

  --r_7 master_run cascaded wait assignment, which is an e_assign
  r_7 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 OR NOT pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 OR NOT pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 OR NOT pixel_buffer_avalon_pixel_buffer_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pixel_buffer_avalon_pixel_buffer_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_master_run <= r_7;
  --optimize select-logic by passing only those address bits which matter.
  internal_pixel_buffer_avalon_pixel_buffer_master_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("000000000") & pixel_buffer_avalon_pixel_buffer_master_address(22 DOWNTO 0));
  --pixel_buffer_avalon_pixel_buffer_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pixel_buffer_avalon_pixel_buffer_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pixel_buffer_avalon_pixel_buffer_master_read_but_no_slave_selected <= (pixel_buffer_avalon_pixel_buffer_master_read AND pixel_buffer_avalon_pixel_buffer_master_run) AND NOT pixel_buffer_avalon_pixel_buffer_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_master_is_granted_some_slave <= pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pixel_buffer_avalon_pixel_buffer_master_readdatavalid <= pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_master_readdatavalid <= pixel_buffer_avalon_pixel_buffer_master_read_but_no_slave_selected OR pre_flush_pixel_buffer_avalon_pixel_buffer_master_readdatavalid;
  --pixel_buffer/avalon_pixel_buffer_master readdata mux, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_master_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_pixel_buffer_avalon_pixel_buffer_master_waitrequest <= NOT pixel_buffer_avalon_pixel_buffer_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pixel_buffer_avalon_pixel_buffer_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_pixel_buffer_avalon_pixel_buffer_master_latency_counter <= p1_pixel_buffer_avalon_pixel_buffer_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pixel_buffer_avalon_pixel_buffer_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((pixel_buffer_avalon_pixel_buffer_master_run AND pixel_buffer_avalon_pixel_buffer_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_pixel_buffer_avalon_pixel_buffer_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_pixel_buffer_avalon_pixel_buffer_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  pixel_buffer_avalon_pixel_buffer_master_address_to_slave <= internal_pixel_buffer_avalon_pixel_buffer_master_address_to_slave;
  --vhdl renameroo for output signals
  pixel_buffer_avalon_pixel_buffer_master_latency_counter <= internal_pixel_buffer_avalon_pixel_buffer_master_latency_counter;
  --vhdl renameroo for output signals
  pixel_buffer_avalon_pixel_buffer_master_waitrequest <= internal_pixel_buffer_avalon_pixel_buffer_master_waitrequest;
--synthesis translate_off
    --pixel_buffer_avalon_pixel_buffer_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pixel_buffer_avalon_pixel_buffer_master_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pixel_buffer_avalon_pixel_buffer_master_address_last_time <= pixel_buffer_avalon_pixel_buffer_master_address;
      end if;

    end process;

    --pixel_buffer/avalon_pixel_buffer_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pixel_buffer_avalon_pixel_buffer_master_waitrequest AND (pixel_buffer_avalon_pixel_buffer_master_read);
      end if;

    end process;

    --pixel_buffer_avalon_pixel_buffer_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pixel_buffer_avalon_pixel_buffer_master_address /= pixel_buffer_avalon_pixel_buffer_master_address_last_time))))) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("pixel_buffer_avalon_pixel_buffer_master_address did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pixel_buffer_avalon_pixel_buffer_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pixel_buffer_avalon_pixel_buffer_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pixel_buffer_avalon_pixel_buffer_master_read_last_time <= pixel_buffer_avalon_pixel_buffer_master_read;
      end if;

    end process;

    --pixel_buffer_avalon_pixel_buffer_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pixel_buffer_avalon_pixel_buffer_master_read) /= std_logic'(pixel_buffer_avalon_pixel_buffer_master_read_last_time)))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("pixel_buffer_avalon_pixel_buffer_master_read did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pixel_buffer_avalon_pixel_buffer_source_arbitrator is 
        port (
              -- inputs:
                 signal alpha_blending_avalon_background_sink_ready_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_source_endofpacket : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_source_startofpacket : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_source_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pixel_buffer_avalon_pixel_buffer_source_ready : OUT STD_LOGIC
              );
end entity pixel_buffer_avalon_pixel_buffer_source_arbitrator;


architecture europa of pixel_buffer_avalon_pixel_buffer_source_arbitrator is

begin

  --mux pixel_buffer_avalon_pixel_buffer_source_ready, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_source_ready <= alpha_blending_avalon_background_sink_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ps2_avalon_ps2_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ps2_avalon_ps2_slave_irq : IN STD_LOGIC;
                 signal ps2_avalon_ps2_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ps2_avalon_ps2_slave_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                 signal d1_ps2_avalon_ps2_slave_end_xfer : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_address : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ps2_avalon_ps2_slave_chipselect : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_irq_from_sa : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_read : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ps2_avalon_ps2_slave_reset : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_write : OUT STD_LOGIC;
                 signal ps2_avalon_ps2_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : OUT STD_LOGIC
              );
end entity ps2_avalon_ps2_slave_arbitrator;


architecture europa of ps2_avalon_ps2_slave_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal internal_ps2_avalon_ps2_slave_waitrequest_from_sa :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_allgrants :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_any_continuerequest :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_arb_counter_enable :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ps2_avalon_ps2_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ps2_avalon_ps2_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ps2_avalon_ps2_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_begins_xfer :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_end_xfer :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_firsttransfer :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_grant_vector :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_in_a_read_cycle :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_in_a_write_cycle :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_master_qreq_vector :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_non_bursting_master_requests :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_reg_firsttransfer :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_slavearbiterlockenable :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_unreg_firsttransfer :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_waits_for_read :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_ps2_avalon_ps2_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal wait_for_ps2_avalon_ps2_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ps2_avalon_ps2_slave_end_xfer;
    end if;

  end process;

  ps2_avalon_ps2_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_ps2_avalon_ps2_slave);
  --assign ps2_avalon_ps2_slave_readdata_from_sa = ps2_avalon_ps2_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  ps2_avalon_ps2_slave_readdata_from_sa <= ps2_avalon_ps2_slave_readdata;
  internal_cpu_data_master_requests_ps2_avalon_ps2_slave <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("110100000011000111110000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign ps2_avalon_ps2_slave_waitrequest_from_sa = ps2_avalon_ps2_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_ps2_avalon_ps2_slave_waitrequest_from_sa <= ps2_avalon_ps2_slave_waitrequest;
  --registered rdv signal_name registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave assignment, which is an e_assign
  registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave <= cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register_in;
  --ps2_avalon_ps2_slave_arb_share_counter set values, which is an e_mux
  ps2_avalon_ps2_slave_arb_share_set_values <= std_logic_vector'("001");
  --ps2_avalon_ps2_slave_non_bursting_master_requests mux, which is an e_mux
  ps2_avalon_ps2_slave_non_bursting_master_requests <= internal_cpu_data_master_requests_ps2_avalon_ps2_slave;
  --ps2_avalon_ps2_slave_any_bursting_master_saved_grant mux, which is an e_mux
  ps2_avalon_ps2_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --ps2_avalon_ps2_slave_arb_share_counter_next_value assignment, which is an e_assign
  ps2_avalon_ps2_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(ps2_avalon_ps2_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (ps2_avalon_ps2_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(ps2_avalon_ps2_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (ps2_avalon_ps2_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --ps2_avalon_ps2_slave_allgrants all slave grants, which is an e_mux
  ps2_avalon_ps2_slave_allgrants <= ps2_avalon_ps2_slave_grant_vector;
  --ps2_avalon_ps2_slave_end_xfer assignment, which is an e_assign
  ps2_avalon_ps2_slave_end_xfer <= NOT ((ps2_avalon_ps2_slave_waits_for_read OR ps2_avalon_ps2_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_ps2_avalon_ps2_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ps2_avalon_ps2_slave <= ps2_avalon_ps2_slave_end_xfer AND (((NOT ps2_avalon_ps2_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ps2_avalon_ps2_slave_arb_share_counter arbitration counter enable, which is an e_assign
  ps2_avalon_ps2_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ps2_avalon_ps2_slave AND ps2_avalon_ps2_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_ps2_avalon_ps2_slave AND NOT ps2_avalon_ps2_slave_non_bursting_master_requests));
  --ps2_avalon_ps2_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ps2_avalon_ps2_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(ps2_avalon_ps2_slave_arb_counter_enable) = '1' then 
        ps2_avalon_ps2_slave_arb_share_counter <= ps2_avalon_ps2_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ps2_avalon_ps2_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ps2_avalon_ps2_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((ps2_avalon_ps2_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_ps2_avalon_ps2_slave)) OR ((end_xfer_arb_share_counter_term_ps2_avalon_ps2_slave AND NOT ps2_avalon_ps2_slave_non_bursting_master_requests)))) = '1' then 
        ps2_avalon_ps2_slave_slavearbiterlockenable <= or_reduce(ps2_avalon_ps2_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master ps2/avalon_ps2_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= ps2_avalon_ps2_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --ps2_avalon_ps2_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ps2_avalon_ps2_slave_slavearbiterlockenable2 <= or_reduce(ps2_avalon_ps2_slave_arb_share_counter_next_value);
  --cpu/data_master ps2/avalon_ps2_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= ps2_avalon_ps2_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --ps2_avalon_ps2_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  ps2_avalon_ps2_slave_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_ps2_avalon_ps2_slave <= internal_cpu_data_master_requests_ps2_avalon_ps2_slave AND NOT ((((cpu_data_master_read AND (cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register))) OR (((NOT cpu_data_master_waitrequest) AND cpu_data_master_write))));
  --cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register_in <= ((internal_cpu_data_master_granted_ps2_avalon_ps2_slave AND cpu_data_master_read) AND NOT ps2_avalon_ps2_slave_waits_for_read) AND NOT (cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register);
  --shift register p1 cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register) & A_ToStdLogicVector(cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register_in)));
  --cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register <= p1_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_ps2_avalon_ps2_slave, which is an e_mux
  cpu_data_master_read_data_valid_ps2_avalon_ps2_slave <= cpu_data_master_read_data_valid_ps2_avalon_ps2_slave_shift_register;
  --ps2_avalon_ps2_slave_writedata mux, which is an e_mux
  ps2_avalon_ps2_slave_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_ps2_avalon_ps2_slave <= internal_cpu_data_master_qualified_request_ps2_avalon_ps2_slave;
  --cpu/data_master saved-grant ps2/avalon_ps2_slave, which is an e_assign
  cpu_data_master_saved_grant_ps2_avalon_ps2_slave <= internal_cpu_data_master_requests_ps2_avalon_ps2_slave;
  --allow new arb cycle for ps2/avalon_ps2_slave, which is an e_assign
  ps2_avalon_ps2_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  ps2_avalon_ps2_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  ps2_avalon_ps2_slave_master_qreq_vector <= std_logic'('1');
  --~ps2_avalon_ps2_slave_reset assignment, which is an e_assign
  ps2_avalon_ps2_slave_reset <= NOT reset_n;
  ps2_avalon_ps2_slave_chipselect <= internal_cpu_data_master_granted_ps2_avalon_ps2_slave;
  --ps2_avalon_ps2_slave_firsttransfer first transaction, which is an e_assign
  ps2_avalon_ps2_slave_firsttransfer <= A_WE_StdLogic((std_logic'(ps2_avalon_ps2_slave_begins_xfer) = '1'), ps2_avalon_ps2_slave_unreg_firsttransfer, ps2_avalon_ps2_slave_reg_firsttransfer);
  --ps2_avalon_ps2_slave_unreg_firsttransfer first transaction, which is an e_assign
  ps2_avalon_ps2_slave_unreg_firsttransfer <= NOT ((ps2_avalon_ps2_slave_slavearbiterlockenable AND ps2_avalon_ps2_slave_any_continuerequest));
  --ps2_avalon_ps2_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ps2_avalon_ps2_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ps2_avalon_ps2_slave_begins_xfer) = '1' then 
        ps2_avalon_ps2_slave_reg_firsttransfer <= ps2_avalon_ps2_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ps2_avalon_ps2_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ps2_avalon_ps2_slave_beginbursttransfer_internal <= ps2_avalon_ps2_slave_begins_xfer;
  --ps2_avalon_ps2_slave_read assignment, which is an e_mux
  ps2_avalon_ps2_slave_read <= internal_cpu_data_master_granted_ps2_avalon_ps2_slave AND cpu_data_master_read;
  --ps2_avalon_ps2_slave_write assignment, which is an e_mux
  ps2_avalon_ps2_slave_write <= internal_cpu_data_master_granted_ps2_avalon_ps2_slave AND cpu_data_master_write;
  shifted_address_to_ps2_avalon_ps2_slave_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --ps2_avalon_ps2_slave_address mux, which is an e_mux
  ps2_avalon_ps2_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_ps2_avalon_ps2_slave_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_ps2_avalon_ps2_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ps2_avalon_ps2_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ps2_avalon_ps2_slave_end_xfer <= ps2_avalon_ps2_slave_end_xfer;
    end if;

  end process;

  --ps2_avalon_ps2_slave_waits_for_read in a cycle, which is an e_mux
  ps2_avalon_ps2_slave_waits_for_read <= ps2_avalon_ps2_slave_in_a_read_cycle AND internal_ps2_avalon_ps2_slave_waitrequest_from_sa;
  --ps2_avalon_ps2_slave_in_a_read_cycle assignment, which is an e_assign
  ps2_avalon_ps2_slave_in_a_read_cycle <= internal_cpu_data_master_granted_ps2_avalon_ps2_slave AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ps2_avalon_ps2_slave_in_a_read_cycle;
  --ps2_avalon_ps2_slave_waits_for_write in a cycle, which is an e_mux
  ps2_avalon_ps2_slave_waits_for_write <= ps2_avalon_ps2_slave_in_a_write_cycle AND internal_ps2_avalon_ps2_slave_waitrequest_from_sa;
  --ps2_avalon_ps2_slave_in_a_write_cycle assignment, which is an e_assign
  ps2_avalon_ps2_slave_in_a_write_cycle <= internal_cpu_data_master_granted_ps2_avalon_ps2_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ps2_avalon_ps2_slave_in_a_write_cycle;
  wait_for_ps2_avalon_ps2_slave_counter <= std_logic'('0');
  --ps2_avalon_ps2_slave_byteenable byte enable port mux, which is an e_mux
  ps2_avalon_ps2_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ps2_avalon_ps2_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --assign ps2_avalon_ps2_slave_irq_from_sa = ps2_avalon_ps2_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  ps2_avalon_ps2_slave_irq_from_sa <= ps2_avalon_ps2_slave_irq;
  --vhdl renameroo for output signals
  cpu_data_master_granted_ps2_avalon_ps2_slave <= internal_cpu_data_master_granted_ps2_avalon_ps2_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_ps2_avalon_ps2_slave <= internal_cpu_data_master_qualified_request_ps2_avalon_ps2_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_ps2_avalon_ps2_slave <= internal_cpu_data_master_requests_ps2_avalon_ps2_slave;
  --vhdl renameroo for output signals
  ps2_avalon_ps2_slave_waitrequest_from_sa <= internal_ps2_avalon_ps2_slave_waitrequest_from_sa;
--synthesis translate_off
    --ps2/avalon_ps2_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_sdram_s1_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1_module;


architecture europa of rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1_module;


architecture europa of rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sdram_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal membuffer_0_avalon_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal membuffer_0_avalon_master_read : IN STD_LOGIC;
                 signal membuffer_0_avalon_master_write : IN STD_LOGIC;
                 signal membuffer_0_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal membuffer_0_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pixel_buffer_avalon_pixel_buffer_master_arbiterlock : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_latency_counter : IN STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_readdatavalid : IN STD_LOGIC;
                 signal sdram_s1_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_byteenable_sdram_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_granted_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_sdram_s1 : OUT STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                 signal membuffer_0_byteenable_sdram_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal membuffer_0_granted_sdram_s1 : OUT STD_LOGIC;
                 signal membuffer_0_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal membuffer_0_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal membuffer_0_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal membuffer_0_requests_sdram_s1 : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 : OUT STD_LOGIC;
                 signal sdram_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal sdram_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sdram_s1_chipselect : OUT STD_LOGIC;
                 signal sdram_s1_read_n : OUT STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sdram_s1_reset_n : OUT STD_LOGIC;
                 signal sdram_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal sdram_s1_write_n : OUT STD_LOGIC;
                 signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sdram_s1_arbitrator;


architecture europa of sdram_s1_arbitrator is
component rdv_fifo_for_cpu_data_master_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_sdram_s1_module;

component rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1_module;

component rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_sdram_s1_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_byteenable_sdram_s1_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal cpu_data_master_saved_grant_sdram_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sdram_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_byteenable_sdram_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_data_master_granted_sdram_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal internal_cpu_data_master_requests_sdram_s1 :  STD_LOGIC;
                signal internal_membuffer_0_byteenable_sdram_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_membuffer_0_granted_sdram_s1 :  STD_LOGIC;
                signal internal_membuffer_0_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_membuffer_0_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal internal_membuffer_0_requests_sdram_s1 :  STD_LOGIC;
                signal internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 :  STD_LOGIC;
                signal internal_pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 :  STD_LOGIC;
                signal internal_sdram_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_cpu_data_master_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_membuffer_0_avalon_master_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_pixel_buffer_avalon_pixel_buffer_master_granted_slave_sdram_s1 :  STD_LOGIC;
                signal membuffer_0_avalon_master_arbiterlock :  STD_LOGIC;
                signal membuffer_0_avalon_master_arbiterlock2 :  STD_LOGIC;
                signal membuffer_0_avalon_master_continuerequest :  STD_LOGIC;
                signal membuffer_0_byteenable_sdram_s1_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal membuffer_0_byteenable_sdram_s1_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal membuffer_0_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal membuffer_0_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal membuffer_0_saved_grant_sdram_s1 :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_arbiterlock2 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_continuerequest :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_saved_grant_sdram_s1 :  STD_LOGIC;
                signal saved_chosen_master_btw_pixel_buffer_avalon_pixel_buffer_master_and_sdram_s1 :  STD_LOGIC;
                signal sdram_s1_allgrants :  STD_LOGIC;
                signal sdram_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sdram_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sdram_s1_any_continuerequest :  STD_LOGIC;
                signal sdram_s1_arb_addend :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_arb_counter_enable :  STD_LOGIC;
                signal sdram_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_arb_winner :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal sdram_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sdram_s1_begins_xfer :  STD_LOGIC;
                signal sdram_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal sdram_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_end_xfer :  STD_LOGIC;
                signal sdram_s1_firsttransfer :  STD_LOGIC;
                signal sdram_s1_grant_vector :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_in_a_read_cycle :  STD_LOGIC;
                signal sdram_s1_in_a_write_cycle :  STD_LOGIC;
                signal sdram_s1_master_qreq_vector :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal sdram_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sdram_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal sdram_s1_reg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sdram_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sdram_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sdram_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_waits_for_read :  STD_LOGIC;
                signal sdram_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sdram_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_membuffer_0_avalon_master :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_pixel_buffer_avalon_pixel_buffer_master :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal wait_for_sdram_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sdram_s1_end_xfer;
    end if;

  end process;

  sdram_s1_begins_xfer <= NOT d1_reasons_to_wait AND (((internal_cpu_data_master_qualified_request_sdram_s1 OR internal_membuffer_0_qualified_request_sdram_s1) OR internal_pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1));
  --assign sdram_s1_readdata_from_sa = sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdata_from_sa <= sdram_s1_readdata;
  internal_cpu_data_master_requests_sdram_s1 <= to_std_logic(((Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_address_to_slave(23)) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("000000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign sdram_s1_waitrequest_from_sa = sdram_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_sdram_s1_waitrequest_from_sa <= sdram_s1_waitrequest;
  --assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdatavalid_from_sa <= sdram_s1_readdatavalid;
  --sdram_s1_arb_share_counter set values, which is an e_mux
  sdram_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_membuffer_0_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_membuffer_0_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_membuffer_0_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001"))))))), 3);
  --sdram_s1_non_bursting_master_requests mux, which is an e_mux
  sdram_s1_non_bursting_master_requests <= (((((((internal_cpu_data_master_requests_sdram_s1 OR internal_membuffer_0_requests_sdram_s1) OR internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1) OR internal_cpu_data_master_requests_sdram_s1) OR internal_membuffer_0_requests_sdram_s1) OR internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1) OR internal_cpu_data_master_requests_sdram_s1) OR internal_membuffer_0_requests_sdram_s1) OR internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1;
  --sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sdram_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  sdram_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sdram_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sdram_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sdram_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --sdram_s1_allgrants all slave grants, which is an e_mux
  sdram_s1_allgrants <= ((((((((or_reduce(sdram_s1_grant_vector)) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector));
  --sdram_s1_end_xfer assignment, which is an e_assign
  sdram_s1_end_xfer <= NOT ((sdram_s1_waits_for_read OR sdram_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sdram_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sdram_s1 <= sdram_s1_end_xfer AND (((NOT sdram_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sdram_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sdram_s1 AND sdram_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests));
  --sdram_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_arb_counter_enable) = '1' then 
        sdram_s1_arb_share_counter <= sdram_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sdram_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_sdram_s1)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests)))) = '1' then 
        sdram_s1_slavearbiterlockenable <= or_reduce(sdram_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master sdram/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= sdram_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sdram_s1_slavearbiterlockenable2 <= or_reduce(sdram_s1_arb_share_counter_next_value);
  --cpu/data_master sdram/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --membuffer_0/avalon_master sdram/s1 arbiterlock, which is an e_assign
  membuffer_0_avalon_master_arbiterlock <= sdram_s1_slavearbiterlockenable AND membuffer_0_avalon_master_continuerequest;
  --membuffer_0/avalon_master sdram/s1 arbiterlock2, which is an e_assign
  membuffer_0_avalon_master_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND membuffer_0_avalon_master_continuerequest;
  --membuffer_0/avalon_master granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_membuffer_0_avalon_master_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_membuffer_0_avalon_master_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(membuffer_0_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_membuffer_0_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_membuffer_0_avalon_master_granted_slave_sdram_s1))))));
    end if;

  end process;

  --membuffer_0_avalon_master_continuerequest continued request, which is an e_mux
  membuffer_0_avalon_master_continuerequest <= ((last_cycle_membuffer_0_avalon_master_granted_slave_sdram_s1 AND internal_membuffer_0_requests_sdram_s1)) OR ((last_cycle_membuffer_0_avalon_master_granted_slave_sdram_s1 AND internal_membuffer_0_requests_sdram_s1));
  --sdram_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  sdram_s1_any_continuerequest <= ((((membuffer_0_avalon_master_continuerequest OR pixel_buffer_avalon_pixel_buffer_master_continuerequest) OR cpu_data_master_continuerequest) OR pixel_buffer_avalon_pixel_buffer_master_continuerequest) OR cpu_data_master_continuerequest) OR membuffer_0_avalon_master_continuerequest;
  --pixel_buffer/avalon_pixel_buffer_master sdram/s1 arbiterlock2, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_master_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND pixel_buffer_avalon_pixel_buffer_master_continuerequest;
  --pixel_buffer/avalon_pixel_buffer_master granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pixel_buffer_avalon_pixel_buffer_master_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pixel_buffer_avalon_pixel_buffer_master_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pixel_buffer_avalon_pixel_buffer_master_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pixel_buffer_avalon_pixel_buffer_master_granted_slave_sdram_s1))))));
    end if;

  end process;

  --pixel_buffer_avalon_pixel_buffer_master_continuerequest continued request, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_master_continuerequest <= ((last_cycle_pixel_buffer_avalon_pixel_buffer_master_granted_slave_sdram_s1 AND internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1)) OR ((last_cycle_pixel_buffer_avalon_pixel_buffer_master_granted_slave_sdram_s1 AND internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1));
  internal_cpu_data_master_qualified_request_sdram_s1 <= internal_cpu_data_master_requests_sdram_s1 AND NOT ((((((cpu_data_master_read AND ((NOT cpu_data_master_waitrequest OR (internal_cpu_data_master_read_data_valid_sdram_s1_shift_register))))) OR (((((NOT cpu_data_master_waitrequest OR cpu_data_master_no_byte_enables_and_last_term) OR NOT(or_reduce(internal_cpu_data_master_byteenable_sdram_s1)))) AND cpu_data_master_write))) OR membuffer_0_avalon_master_arbiterlock) OR ((pixel_buffer_avalon_pixel_buffer_master_arbiterlock AND (saved_chosen_master_btw_pixel_buffer_avalon_pixel_buffer_master_and_sdram_s1)))));
  --unique name for sdram_s1_move_on_to_next_transaction, which is an e_assign
  sdram_s1_move_on_to_next_transaction <= sdram_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_sdram_s1 : rdv_fifo_for_cpu_data_master_to_sdram_s1_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => internal_cpu_data_master_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  internal_cpu_data_master_read_data_valid_sdram_s1_shift_register <= NOT cpu_data_master_rdv_fifo_empty_sdram_s1;
  --local readdatavalid cpu_data_master_read_data_valid_sdram_s1, which is an e_mux
  cpu_data_master_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND cpu_data_master_rdv_fifo_output_from_sdram_s1)) AND NOT cpu_data_master_rdv_fifo_empty_sdram_s1;
  --sdram_s1_writedata mux, which is an e_mux
  sdram_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sdram_s1)) = '1'), cpu_data_master_dbs_write_16, membuffer_0_dbs_write_16);
  internal_membuffer_0_requests_sdram_s1 <= to_std_logic(((Std_Logic_Vector'(membuffer_0_avalon_master_address_to_slave(31 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND ((membuffer_0_avalon_master_read OR membuffer_0_avalon_master_write));
  --cpu/data_master granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_data_master_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_data_master_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_data_master_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_cpu_data_master_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_data_master_granted_slave_sdram_s1))))));
    end if;

  end process;

  --cpu_data_master_continuerequest continued request, which is an e_mux
  cpu_data_master_continuerequest <= ((last_cycle_cpu_data_master_granted_slave_sdram_s1 AND internal_cpu_data_master_requests_sdram_s1)) OR ((last_cycle_cpu_data_master_granted_slave_sdram_s1 AND internal_cpu_data_master_requests_sdram_s1));
  internal_membuffer_0_qualified_request_sdram_s1 <= internal_membuffer_0_requests_sdram_s1 AND NOT (((((membuffer_0_avalon_master_read AND (internal_membuffer_0_read_data_valid_sdram_s1_shift_register))) OR cpu_data_master_arbiterlock) OR ((pixel_buffer_avalon_pixel_buffer_master_arbiterlock AND (saved_chosen_master_btw_pixel_buffer_avalon_pixel_buffer_master_and_sdram_s1)))));
  --rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1 : rdv_fifo_for_membuffer_0_avalon_master_to_sdram_s1_module
    port map(
      data_out => membuffer_0_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => membuffer_0_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_membuffer_0_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  internal_membuffer_0_read_data_valid_sdram_s1_shift_register <= NOT membuffer_0_rdv_fifo_empty_sdram_s1;
  --local readdatavalid membuffer_0_read_data_valid_sdram_s1, which is an e_mux
  membuffer_0_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND membuffer_0_rdv_fifo_output_from_sdram_s1)) AND NOT membuffer_0_rdv_fifo_empty_sdram_s1;
  internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 <= ((to_std_logic(((Std_Logic_Vector'(pixel_buffer_avalon_pixel_buffer_master_address_to_slave(31 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (pixel_buffer_avalon_pixel_buffer_master_read))) AND pixel_buffer_avalon_pixel_buffer_master_read;
  internal_pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 <= internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 AND NOT (((((pixel_buffer_avalon_pixel_buffer_master_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pixel_buffer_avalon_pixel_buffer_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pixel_buffer_avalon_pixel_buffer_master_latency_counter)))))))))) OR cpu_data_master_arbiterlock) OR membuffer_0_avalon_master_arbiterlock));
  --rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1 : rdv_fifo_for_pixel_buffer_avalon_pixel_buffer_master_to_sdram_s1_module
    port map(
      data_out => pixel_buffer_avalon_pixel_buffer_master_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => pixel_buffer_avalon_pixel_buffer_master_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register <= NOT pixel_buffer_avalon_pixel_buffer_master_rdv_fifo_empty_sdram_s1;
  --local readdatavalid pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1, which is an e_mux
  pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND pixel_buffer_avalon_pixel_buffer_master_rdv_fifo_output_from_sdram_s1)) AND NOT pixel_buffer_avalon_pixel_buffer_master_rdv_fifo_empty_sdram_s1;
  --allow new arb cycle for sdram/s1, which is an e_assign
  sdram_s1_allow_new_arb_cycle <= (NOT cpu_data_master_arbiterlock AND NOT membuffer_0_avalon_master_arbiterlock) AND NOT ((pixel_buffer_avalon_pixel_buffer_master_arbiterlock AND (saved_chosen_master_btw_pixel_buffer_avalon_pixel_buffer_master_and_sdram_s1)));
  --pixel_buffer/avalon_pixel_buffer_master assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(0) <= internal_pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1;
  --pixel_buffer/avalon_pixel_buffer_master grant sdram/s1, which is an e_assign
  internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 <= sdram_s1_grant_vector(0);
  --pixel_buffer/avalon_pixel_buffer_master saved-grant sdram/s1, which is an e_assign
  pixel_buffer_avalon_pixel_buffer_master_saved_grant_sdram_s1 <= sdram_s1_arb_winner(0) AND internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1;
  --saved chosen master btw pixel_buffer/avalon_pixel_buffer_master and sdram/s1, which is an e_assign
  saved_chosen_master_btw_pixel_buffer_avalon_pixel_buffer_master_and_sdram_s1 <= sdram_s1_saved_chosen_master_vector(0);
  --membuffer_0/avalon_master assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(1) <= internal_membuffer_0_qualified_request_sdram_s1;
  --membuffer_0/avalon_master grant sdram/s1, which is an e_assign
  internal_membuffer_0_granted_sdram_s1 <= sdram_s1_grant_vector(1);
  --membuffer_0/avalon_master saved-grant sdram/s1, which is an e_assign
  membuffer_0_saved_grant_sdram_s1 <= sdram_s1_arb_winner(1) AND internal_membuffer_0_requests_sdram_s1;
  --cpu/data_master assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(2) <= internal_cpu_data_master_qualified_request_sdram_s1;
  --cpu/data_master grant sdram/s1, which is an e_assign
  internal_cpu_data_master_granted_sdram_s1 <= sdram_s1_grant_vector(2);
  --cpu/data_master saved-grant sdram/s1, which is an e_assign
  cpu_data_master_saved_grant_sdram_s1 <= sdram_s1_arb_winner(2) AND internal_cpu_data_master_requests_sdram_s1;
  --sdram/s1 chosen-master double-vector, which is an e_assign
  sdram_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sdram_s1_master_qreq_vector & sdram_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sdram_s1_master_qreq_vector & NOT sdram_s1_master_qreq_vector))) + (std_logic_vector'("0000") & (sdram_s1_arb_addend))))), 6);
  --stable onehot encoding of arb winner
  sdram_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((sdram_s1_allow_new_arb_cycle AND or_reduce(sdram_s1_grant_vector)))) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
  --saved sdram_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_saved_chosen_master_vector <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_allow_new_arb_cycle) = '1' then 
        sdram_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_grant_vector)) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sdram_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(2) OR sdram_s1_chosen_master_double_vector(5)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(1) OR sdram_s1_chosen_master_double_vector(4)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(0) OR sdram_s1_chosen_master_double_vector(3)))));
  --sdram/s1 chosen master rotated left, which is an e_assign
  sdram_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("000")), (std_logic_vector'("00000000000000000000000000000") & ((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 3);
  --sdram/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_addend <= std_logic_vector'("001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sdram_s1_grant_vector)) = '1' then 
        sdram_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(sdram_s1_end_xfer) = '1'), sdram_s1_chosen_master_rot_left, sdram_s1_grant_vector);
      end if;
    end if;

  end process;

  --sdram_s1_reset_n assignment, which is an e_assign
  sdram_s1_reset_n <= reset_n;
  sdram_s1_chipselect <= (internal_cpu_data_master_granted_sdram_s1 OR internal_membuffer_0_granted_sdram_s1) OR internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1;
  --sdram_s1_firsttransfer first transaction, which is an e_assign
  sdram_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sdram_s1_begins_xfer) = '1'), sdram_s1_unreg_firsttransfer, sdram_s1_reg_firsttransfer);
  --sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  sdram_s1_unreg_firsttransfer <= NOT ((sdram_s1_slavearbiterlockenable AND sdram_s1_any_continuerequest));
  --sdram_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_begins_xfer) = '1' then 
        sdram_s1_reg_firsttransfer <= sdram_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sdram_s1_beginbursttransfer_internal <= sdram_s1_begins_xfer;
  --sdram_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sdram_s1_arbitration_holdoff_internal <= sdram_s1_begins_xfer AND sdram_s1_firsttransfer;
  --~sdram_s1_read_n assignment, which is an e_mux
  sdram_s1_read_n <= NOT (((((internal_cpu_data_master_granted_sdram_s1 AND cpu_data_master_read)) OR ((internal_membuffer_0_granted_sdram_s1 AND membuffer_0_avalon_master_read))) OR ((internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 AND pixel_buffer_avalon_pixel_buffer_master_read))));
  --~sdram_s1_write_n assignment, which is an e_mux
  sdram_s1_write_n <= NOT ((((internal_cpu_data_master_granted_sdram_s1 AND cpu_data_master_write)) OR ((internal_membuffer_0_granted_sdram_s1 AND membuffer_0_avalon_master_write))));
  shifted_address_to_sdram_s1_from_cpu_data_master <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 24);
  --sdram_s1_address mux, which is an e_mux
  sdram_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sdram_s1)) = '1'), (std_logic_vector'("00000000") & ((A_SRL(shifted_address_to_sdram_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000001"))))), A_WE_StdLogicVector((std_logic'((internal_membuffer_0_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_membuffer_0_avalon_master,std_logic_vector'("00000000000000000000000000000001"))), (A_SRL(shifted_address_to_sdram_s1_from_pixel_buffer_avalon_pixel_buffer_master,std_logic_vector'("00000000000000000000000000000001"))))), 22);
  shifted_address_to_sdram_s1_from_membuffer_0_avalon_master <= A_EXT (Std_Logic_Vector'(A_SRL(membuffer_0_avalon_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(membuffer_0_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 32);
  shifted_address_to_sdram_s1_from_pixel_buffer_avalon_pixel_buffer_master <= pixel_buffer_avalon_pixel_buffer_master_address_to_slave;
  --d1_sdram_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sdram_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sdram_s1_end_xfer <= sdram_s1_end_xfer;
    end if;

  end process;

  --sdram_s1_waits_for_read in a cycle, which is an e_mux
  sdram_s1_waits_for_read <= sdram_s1_in_a_read_cycle AND internal_sdram_s1_waitrequest_from_sa;
  --sdram_s1_in_a_read_cycle assignment, which is an e_assign
  sdram_s1_in_a_read_cycle <= (((internal_cpu_data_master_granted_sdram_s1 AND cpu_data_master_read)) OR ((internal_membuffer_0_granted_sdram_s1 AND membuffer_0_avalon_master_read))) OR ((internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 AND pixel_buffer_avalon_pixel_buffer_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sdram_s1_in_a_read_cycle;
  --sdram_s1_waits_for_write in a cycle, which is an e_mux
  sdram_s1_waits_for_write <= sdram_s1_in_a_write_cycle AND internal_sdram_s1_waitrequest_from_sa;
  --sdram_s1_in_a_write_cycle assignment, which is an e_assign
  sdram_s1_in_a_write_cycle <= ((internal_cpu_data_master_granted_sdram_s1 AND cpu_data_master_write)) OR ((internal_membuffer_0_granted_sdram_s1 AND membuffer_0_avalon_master_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sdram_s1_in_a_write_cycle;
  wait_for_sdram_s1_counter <= std_logic'('0');
  --~sdram_s1_byteenable_n byte enable port mux, which is an e_mux
  sdram_s1_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_byteenable_sdram_s1)), A_WE_StdLogicVector((std_logic'((internal_membuffer_0_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_membuffer_0_byteenable_sdram_s1)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))), 2);
  (cpu_data_master_byteenable_sdram_s1_segment_1(1), cpu_data_master_byteenable_sdram_s1_segment_1(0), cpu_data_master_byteenable_sdram_s1_segment_0(1), cpu_data_master_byteenable_sdram_s1_segment_0(0)) <= cpu_data_master_byteenable;
  internal_cpu_data_master_byteenable_sdram_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_byteenable_sdram_s1_segment_0, cpu_data_master_byteenable_sdram_s1_segment_1);
  (membuffer_0_byteenable_sdram_s1_segment_1(1), membuffer_0_byteenable_sdram_s1_segment_1(0), membuffer_0_byteenable_sdram_s1_segment_0(1), membuffer_0_byteenable_sdram_s1_segment_0(0)) <= A_REP(std_logic'('1'), 4);
  internal_membuffer_0_byteenable_sdram_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(membuffer_0_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), membuffer_0_byteenable_sdram_s1_segment_0, membuffer_0_byteenable_sdram_s1_segment_1);
  --vhdl renameroo for output signals
  cpu_data_master_byteenable_sdram_s1 <= internal_cpu_data_master_byteenable_sdram_s1;
  --vhdl renameroo for output signals
  cpu_data_master_granted_sdram_s1 <= internal_cpu_data_master_granted_sdram_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_sdram_s1 <= internal_cpu_data_master_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  cpu_data_master_read_data_valid_sdram_s1_shift_register <= internal_cpu_data_master_read_data_valid_sdram_s1_shift_register;
  --vhdl renameroo for output signals
  cpu_data_master_requests_sdram_s1 <= internal_cpu_data_master_requests_sdram_s1;
  --vhdl renameroo for output signals
  membuffer_0_byteenable_sdram_s1 <= internal_membuffer_0_byteenable_sdram_s1;
  --vhdl renameroo for output signals
  membuffer_0_granted_sdram_s1 <= internal_membuffer_0_granted_sdram_s1;
  --vhdl renameroo for output signals
  membuffer_0_qualified_request_sdram_s1 <= internal_membuffer_0_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  membuffer_0_read_data_valid_sdram_s1_shift_register <= internal_membuffer_0_read_data_valid_sdram_s1_shift_register;
  --vhdl renameroo for output signals
  membuffer_0_requests_sdram_s1 <= internal_membuffer_0_requests_sdram_s1;
  --vhdl renameroo for output signals
  pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 <= internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1;
  --vhdl renameroo for output signals
  pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 <= internal_pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 <= internal_pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1;
  --vhdl renameroo for output signals
  sdram_s1_waitrequest_from_sa <= internal_sdram_s1_waitrequest_from_sa;
--synthesis translate_off
    --sdram/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("00000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_granted_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_membuffer_0_granted_sdram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("00000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_data_master_saved_grant_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(membuffer_0_saved_grant_sdram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(pixel_buffer_avalon_pixel_buffer_master_saved_grant_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sram_avalon_sram_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sram_avalon_sram_slave_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal cpu_data_master_byteenable_sram_avalon_sram_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cpu_data_master_granted_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal cpu_data_master_requests_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal cpu_instruction_master_granted_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal d1_sram_avalon_sram_slave_end_xfer : OUT STD_LOGIC;
                 signal registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave : OUT STD_LOGIC;
                 signal sram_avalon_sram_slave_address : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal sram_avalon_sram_slave_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sram_avalon_sram_slave_read : OUT STD_LOGIC;
                 signal sram_avalon_sram_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sram_avalon_sram_slave_reset : OUT STD_LOGIC;
                 signal sram_avalon_sram_slave_write : OUT STD_LOGIC;
                 signal sram_avalon_sram_slave_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sram_avalon_sram_slave_arbitrator;


architecture europa of sram_avalon_sram_slave_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_byteenable_sram_avalon_sram_slave_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_byteenable_sram_avalon_sram_slave_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register_in :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_sram_avalon_sram_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sram_avalon_sram_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_byteenable_sram_avalon_sram_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_cpu_data_master_granted_sram_avalon_sram_slave :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_sram_avalon_sram_slave :  STD_LOGIC;
                signal internal_cpu_data_master_requests_sram_avalon_sram_slave :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_sram_avalon_sram_slave :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_sram_avalon_sram_slave :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_sram_avalon_sram_slave :  STD_LOGIC;
                signal last_cycle_cpu_data_master_granted_slave_sram_avalon_sram_slave :  STD_LOGIC;
                signal last_cycle_cpu_instruction_master_granted_slave_sram_avalon_sram_slave :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal shifted_address_to_sram_avalon_sram_slave_from_cpu_data_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal shifted_address_to_sram_avalon_sram_slave_from_cpu_instruction_master :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal sram_avalon_sram_slave_allgrants :  STD_LOGIC;
                signal sram_avalon_sram_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal sram_avalon_sram_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sram_avalon_sram_slave_any_continuerequest :  STD_LOGIC;
                signal sram_avalon_sram_slave_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_avalon_sram_slave_arb_counter_enable :  STD_LOGIC;
                signal sram_avalon_sram_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sram_avalon_sram_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sram_avalon_sram_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sram_avalon_sram_slave_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_avalon_sram_slave_arbitration_holdoff_internal :  STD_LOGIC;
                signal sram_avalon_sram_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal sram_avalon_sram_slave_begins_xfer :  STD_LOGIC;
                signal sram_avalon_sram_slave_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sram_avalon_sram_slave_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_avalon_sram_slave_end_xfer :  STD_LOGIC;
                signal sram_avalon_sram_slave_firsttransfer :  STD_LOGIC;
                signal sram_avalon_sram_slave_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_avalon_sram_slave_in_a_read_cycle :  STD_LOGIC;
                signal sram_avalon_sram_slave_in_a_write_cycle :  STD_LOGIC;
                signal sram_avalon_sram_slave_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_avalon_sram_slave_non_bursting_master_requests :  STD_LOGIC;
                signal sram_avalon_sram_slave_reg_firsttransfer :  STD_LOGIC;
                signal sram_avalon_sram_slave_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_avalon_sram_slave_slavearbiterlockenable :  STD_LOGIC;
                signal sram_avalon_sram_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal sram_avalon_sram_slave_unreg_firsttransfer :  STD_LOGIC;
                signal sram_avalon_sram_slave_waits_for_read :  STD_LOGIC;
                signal sram_avalon_sram_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_sram_avalon_sram_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sram_avalon_sram_slave_end_xfer;
    end if;

  end process;

  sram_avalon_sram_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_data_master_qualified_request_sram_avalon_sram_slave OR internal_cpu_instruction_master_qualified_request_sram_avalon_sram_slave));
  --assign sram_avalon_sram_slave_readdata_from_sa = sram_avalon_sram_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sram_avalon_sram_slave_readdata_from_sa <= sram_avalon_sram_slave_readdata;
  internal_cpu_data_master_requests_sram_avalon_sram_slave <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(23 DOWNTO 19) & std_logic_vector'("0000000000000000000")) = std_logic_vector'("110010000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --registered rdv signal_name registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave assignment, which is an e_assign
  registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave <= cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register(0);
  --sram_avalon_sram_slave_arb_share_counter set values, which is an e_mux
  sram_avalon_sram_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sram_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_sram_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sram_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_sram_avalon_sram_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001"))))), 3);
  --sram_avalon_sram_slave_non_bursting_master_requests mux, which is an e_mux
  sram_avalon_sram_slave_non_bursting_master_requests <= ((internal_cpu_data_master_requests_sram_avalon_sram_slave OR internal_cpu_instruction_master_requests_sram_avalon_sram_slave) OR internal_cpu_data_master_requests_sram_avalon_sram_slave) OR internal_cpu_instruction_master_requests_sram_avalon_sram_slave;
  --sram_avalon_sram_slave_any_bursting_master_saved_grant mux, which is an e_mux
  sram_avalon_sram_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --sram_avalon_sram_slave_arb_share_counter_next_value assignment, which is an e_assign
  sram_avalon_sram_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sram_avalon_sram_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sram_avalon_sram_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sram_avalon_sram_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sram_avalon_sram_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --sram_avalon_sram_slave_allgrants all slave grants, which is an e_mux
  sram_avalon_sram_slave_allgrants <= (((or_reduce(sram_avalon_sram_slave_grant_vector)) OR (or_reduce(sram_avalon_sram_slave_grant_vector))) OR (or_reduce(sram_avalon_sram_slave_grant_vector))) OR (or_reduce(sram_avalon_sram_slave_grant_vector));
  --sram_avalon_sram_slave_end_xfer assignment, which is an e_assign
  sram_avalon_sram_slave_end_xfer <= NOT ((sram_avalon_sram_slave_waits_for_read OR sram_avalon_sram_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_sram_avalon_sram_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sram_avalon_sram_slave <= sram_avalon_sram_slave_end_xfer AND (((NOT sram_avalon_sram_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sram_avalon_sram_slave_arb_share_counter arbitration counter enable, which is an e_assign
  sram_avalon_sram_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sram_avalon_sram_slave AND sram_avalon_sram_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_sram_avalon_sram_slave AND NOT sram_avalon_sram_slave_non_bursting_master_requests));
  --sram_avalon_sram_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_avalon_sram_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(sram_avalon_sram_slave_arb_counter_enable) = '1' then 
        sram_avalon_sram_slave_arb_share_counter <= sram_avalon_sram_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sram_avalon_sram_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_avalon_sram_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sram_avalon_sram_slave_master_qreq_vector) AND end_xfer_arb_share_counter_term_sram_avalon_sram_slave)) OR ((end_xfer_arb_share_counter_term_sram_avalon_sram_slave AND NOT sram_avalon_sram_slave_non_bursting_master_requests)))) = '1' then 
        sram_avalon_sram_slave_slavearbiterlockenable <= or_reduce(sram_avalon_sram_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master sram/avalon_sram_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= sram_avalon_sram_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --sram_avalon_sram_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sram_avalon_sram_slave_slavearbiterlockenable2 <= or_reduce(sram_avalon_sram_slave_arb_share_counter_next_value);
  --cpu/data_master sram/avalon_sram_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= sram_avalon_sram_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --cpu/instruction_master sram/avalon_sram_slave arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= sram_avalon_sram_slave_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master sram/avalon_sram_slave arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= sram_avalon_sram_slave_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master granted sram/avalon_sram_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_instruction_master_granted_slave_sram_avalon_sram_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_instruction_master_granted_slave_sram_avalon_sram_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_instruction_master_saved_grant_sram_avalon_sram_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sram_avalon_sram_slave_arbitration_holdoff_internal OR NOT internal_cpu_instruction_master_requests_sram_avalon_sram_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_instruction_master_granted_slave_sram_avalon_sram_slave))))));
    end if;

  end process;

  --cpu_instruction_master_continuerequest continued request, which is an e_mux
  cpu_instruction_master_continuerequest <= last_cycle_cpu_instruction_master_granted_slave_sram_avalon_sram_slave AND internal_cpu_instruction_master_requests_sram_avalon_sram_slave;
  --sram_avalon_sram_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  sram_avalon_sram_slave_any_continuerequest <= cpu_instruction_master_continuerequest OR cpu_data_master_continuerequest;
  internal_cpu_data_master_qualified_request_sram_avalon_sram_slave <= internal_cpu_data_master_requests_sram_avalon_sram_slave AND NOT (((((cpu_data_master_read AND (or_reduce(cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register)))) OR (((((NOT cpu_data_master_waitrequest OR cpu_data_master_no_byte_enables_and_last_term) OR NOT(or_reduce(internal_cpu_data_master_byteenable_sram_avalon_sram_slave)))) AND cpu_data_master_write))) OR cpu_instruction_master_arbiterlock));
  --cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register_in <= ((internal_cpu_data_master_granted_sram_avalon_sram_slave AND cpu_data_master_read) AND NOT sram_avalon_sram_slave_waits_for_read) AND NOT (or_reduce(cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register));
  --shift register p1 cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register <= A_EXT ((cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register & A_ToStdLogicVector(cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register_in)), 2);
  --cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register <= p1_cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_sram_avalon_sram_slave, which is an e_mux
  cpu_data_master_read_data_valid_sram_avalon_sram_slave <= cpu_data_master_read_data_valid_sram_avalon_sram_slave_shift_register(1);
  --sram_avalon_sram_slave_writedata mux, which is an e_mux
  sram_avalon_sram_slave_writedata <= cpu_data_master_dbs_write_16;
  internal_cpu_instruction_master_requests_sram_avalon_sram_slave <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(23 DOWNTO 19) & std_logic_vector'("0000000000000000000")) = std_logic_vector'("110010000000000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --cpu/data_master granted sram/avalon_sram_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_data_master_granted_slave_sram_avalon_sram_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_data_master_granted_slave_sram_avalon_sram_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_data_master_saved_grant_sram_avalon_sram_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sram_avalon_sram_slave_arbitration_holdoff_internal OR NOT internal_cpu_data_master_requests_sram_avalon_sram_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_data_master_granted_slave_sram_avalon_sram_slave))))));
    end if;

  end process;

  --cpu_data_master_continuerequest continued request, which is an e_mux
  cpu_data_master_continuerequest <= last_cycle_cpu_data_master_granted_slave_sram_avalon_sram_slave AND internal_cpu_data_master_requests_sram_avalon_sram_slave;
  internal_cpu_instruction_master_qualified_request_sram_avalon_sram_slave <= internal_cpu_instruction_master_requests_sram_avalon_sram_slave AND NOT ((((cpu_instruction_master_read AND to_std_logic(((std_logic_vector'("00000000000000000000000000000010")<(std_logic_vector'("000000000000000000000000000000") & (cpu_instruction_master_latency_counter))))))) OR cpu_data_master_arbiterlock));
  --cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register_in <= (internal_cpu_instruction_master_granted_sram_avalon_sram_slave AND cpu_instruction_master_read) AND NOT sram_avalon_sram_slave_waits_for_read;
  --shift register p1 cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register <= A_EXT ((cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register & A_ToStdLogicVector(cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register_in)), 2);
  --cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register <= p1_cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_instruction_master_read_data_valid_sram_avalon_sram_slave, which is an e_mux
  cpu_instruction_master_read_data_valid_sram_avalon_sram_slave <= cpu_instruction_master_read_data_valid_sram_avalon_sram_slave_shift_register(1);
  --allow new arb cycle for sram/avalon_sram_slave, which is an e_assign
  sram_avalon_sram_slave_allow_new_arb_cycle <= NOT cpu_data_master_arbiterlock AND NOT cpu_instruction_master_arbiterlock;
  --cpu/instruction_master assignment into master qualified-requests vector for sram/avalon_sram_slave, which is an e_assign
  sram_avalon_sram_slave_master_qreq_vector(0) <= internal_cpu_instruction_master_qualified_request_sram_avalon_sram_slave;
  --cpu/instruction_master grant sram/avalon_sram_slave, which is an e_assign
  internal_cpu_instruction_master_granted_sram_avalon_sram_slave <= sram_avalon_sram_slave_grant_vector(0);
  --cpu/instruction_master saved-grant sram/avalon_sram_slave, which is an e_assign
  cpu_instruction_master_saved_grant_sram_avalon_sram_slave <= sram_avalon_sram_slave_arb_winner(0) AND internal_cpu_instruction_master_requests_sram_avalon_sram_slave;
  --cpu/data_master assignment into master qualified-requests vector for sram/avalon_sram_slave, which is an e_assign
  sram_avalon_sram_slave_master_qreq_vector(1) <= internal_cpu_data_master_qualified_request_sram_avalon_sram_slave;
  --cpu/data_master grant sram/avalon_sram_slave, which is an e_assign
  internal_cpu_data_master_granted_sram_avalon_sram_slave <= sram_avalon_sram_slave_grant_vector(1);
  --cpu/data_master saved-grant sram/avalon_sram_slave, which is an e_assign
  cpu_data_master_saved_grant_sram_avalon_sram_slave <= sram_avalon_sram_slave_arb_winner(1) AND internal_cpu_data_master_requests_sram_avalon_sram_slave;
  --sram/avalon_sram_slave chosen-master double-vector, which is an e_assign
  sram_avalon_sram_slave_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sram_avalon_sram_slave_master_qreq_vector & sram_avalon_sram_slave_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sram_avalon_sram_slave_master_qreq_vector & NOT sram_avalon_sram_slave_master_qreq_vector))) + (std_logic_vector'("000") & (sram_avalon_sram_slave_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  sram_avalon_sram_slave_arb_winner <= A_WE_StdLogicVector((std_logic'(((sram_avalon_sram_slave_allow_new_arb_cycle AND or_reduce(sram_avalon_sram_slave_grant_vector)))) = '1'), sram_avalon_sram_slave_grant_vector, sram_avalon_sram_slave_saved_chosen_master_vector);
  --saved sram_avalon_sram_slave_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_avalon_sram_slave_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(sram_avalon_sram_slave_allow_new_arb_cycle) = '1' then 
        sram_avalon_sram_slave_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sram_avalon_sram_slave_grant_vector)) = '1'), sram_avalon_sram_slave_grant_vector, sram_avalon_sram_slave_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sram_avalon_sram_slave_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sram_avalon_sram_slave_chosen_master_double_vector(1) OR sram_avalon_sram_slave_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((sram_avalon_sram_slave_chosen_master_double_vector(0) OR sram_avalon_sram_slave_chosen_master_double_vector(2)))));
  --sram/avalon_sram_slave chosen master rotated left, which is an e_assign
  sram_avalon_sram_slave_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sram_avalon_sram_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(sram_avalon_sram_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --sram/avalon_sram_slave's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_avalon_sram_slave_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sram_avalon_sram_slave_grant_vector)) = '1' then 
        sram_avalon_sram_slave_arb_addend <= A_WE_StdLogicVector((std_logic'(sram_avalon_sram_slave_end_xfer) = '1'), sram_avalon_sram_slave_chosen_master_rot_left, sram_avalon_sram_slave_grant_vector);
      end if;
    end if;

  end process;

  --~sram_avalon_sram_slave_reset assignment, which is an e_assign
  sram_avalon_sram_slave_reset <= NOT reset_n;
  --sram_avalon_sram_slave_firsttransfer first transaction, which is an e_assign
  sram_avalon_sram_slave_firsttransfer <= A_WE_StdLogic((std_logic'(sram_avalon_sram_slave_begins_xfer) = '1'), sram_avalon_sram_slave_unreg_firsttransfer, sram_avalon_sram_slave_reg_firsttransfer);
  --sram_avalon_sram_slave_unreg_firsttransfer first transaction, which is an e_assign
  sram_avalon_sram_slave_unreg_firsttransfer <= NOT ((sram_avalon_sram_slave_slavearbiterlockenable AND sram_avalon_sram_slave_any_continuerequest));
  --sram_avalon_sram_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sram_avalon_sram_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sram_avalon_sram_slave_begins_xfer) = '1' then 
        sram_avalon_sram_slave_reg_firsttransfer <= sram_avalon_sram_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sram_avalon_sram_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sram_avalon_sram_slave_beginbursttransfer_internal <= sram_avalon_sram_slave_begins_xfer;
  --sram_avalon_sram_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sram_avalon_sram_slave_arbitration_holdoff_internal <= sram_avalon_sram_slave_begins_xfer AND sram_avalon_sram_slave_firsttransfer;
  --sram_avalon_sram_slave_read assignment, which is an e_mux
  sram_avalon_sram_slave_read <= ((internal_cpu_data_master_granted_sram_avalon_sram_slave AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_sram_avalon_sram_slave AND cpu_instruction_master_read));
  --sram_avalon_sram_slave_write assignment, which is an e_mux
  sram_avalon_sram_slave_write <= internal_cpu_data_master_granted_sram_avalon_sram_slave AND cpu_data_master_write;
  shifted_address_to_sram_avalon_sram_slave_from_cpu_data_master <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 24);
  --sram_avalon_sram_slave_address mux, which is an e_mux
  sram_avalon_sram_slave_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sram_avalon_sram_slave)) = '1'), (A_SRL(shifted_address_to_sram_avalon_sram_slave_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000001"))), (A_SRL(shifted_address_to_sram_avalon_sram_slave_from_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000001")))), 18);
  shifted_address_to_sram_avalon_sram_slave_from_cpu_instruction_master <= A_EXT (Std_Logic_Vector'(A_SRL(cpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(cpu_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 24);
  --d1_sram_avalon_sram_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sram_avalon_sram_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sram_avalon_sram_slave_end_xfer <= sram_avalon_sram_slave_end_xfer;
    end if;

  end process;

  --sram_avalon_sram_slave_waits_for_read in a cycle, which is an e_mux
  sram_avalon_sram_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sram_avalon_sram_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sram_avalon_sram_slave_in_a_read_cycle assignment, which is an e_assign
  sram_avalon_sram_slave_in_a_read_cycle <= ((internal_cpu_data_master_granted_sram_avalon_sram_slave AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_sram_avalon_sram_slave AND cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sram_avalon_sram_slave_in_a_read_cycle;
  --sram_avalon_sram_slave_waits_for_write in a cycle, which is an e_mux
  sram_avalon_sram_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sram_avalon_sram_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sram_avalon_sram_slave_in_a_write_cycle assignment, which is an e_assign
  sram_avalon_sram_slave_in_a_write_cycle <= internal_cpu_data_master_granted_sram_avalon_sram_slave AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sram_avalon_sram_slave_in_a_write_cycle;
  wait_for_sram_avalon_sram_slave_counter <= std_logic'('0');
  --sram_avalon_sram_slave_byteenable byte enable port mux, which is an e_mux
  sram_avalon_sram_slave_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_sram_avalon_sram_slave)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_byteenable_sram_avalon_sram_slave)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  (cpu_data_master_byteenable_sram_avalon_sram_slave_segment_1(1), cpu_data_master_byteenable_sram_avalon_sram_slave_segment_1(0), cpu_data_master_byteenable_sram_avalon_sram_slave_segment_0(1), cpu_data_master_byteenable_sram_avalon_sram_slave_segment_0(0)) <= cpu_data_master_byteenable;
  internal_cpu_data_master_byteenable_sram_avalon_sram_slave <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), cpu_data_master_byteenable_sram_avalon_sram_slave_segment_0, cpu_data_master_byteenable_sram_avalon_sram_slave_segment_1);
  --vhdl renameroo for output signals
  cpu_data_master_byteenable_sram_avalon_sram_slave <= internal_cpu_data_master_byteenable_sram_avalon_sram_slave;
  --vhdl renameroo for output signals
  cpu_data_master_granted_sram_avalon_sram_slave <= internal_cpu_data_master_granted_sram_avalon_sram_slave;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_sram_avalon_sram_slave <= internal_cpu_data_master_qualified_request_sram_avalon_sram_slave;
  --vhdl renameroo for output signals
  cpu_data_master_requests_sram_avalon_sram_slave <= internal_cpu_data_master_requests_sram_avalon_sram_slave;
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_sram_avalon_sram_slave <= internal_cpu_instruction_master_granted_sram_avalon_sram_slave;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_sram_avalon_sram_slave <= internal_cpu_instruction_master_qualified_request_sram_avalon_sram_slave;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_sram_avalon_sram_slave <= internal_cpu_instruction_master_requests_sram_avalon_sram_slave;
--synthesis translate_off
    --sram/avalon_sram_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_granted_sram_avalon_sram_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_instruction_master_granted_sram_avalon_sram_slave))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_data_master_saved_grant_sram_avalon_sram_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_saved_grant_sram_avalon_sram_slave))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity vga_avalon_vga_sink_arbitrator is 
        port (
              -- inputs:
                 signal alpha_blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal alpha_blending_avalon_blended_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal alpha_blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                 signal alpha_blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                 signal alpha_blending_avalon_blended_source_valid : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal vga_avalon_vga_sink_ready : IN STD_LOGIC;

              -- outputs:
                 signal vga_avalon_vga_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                 signal vga_avalon_vga_sink_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal vga_avalon_vga_sink_endofpacket : OUT STD_LOGIC;
                 signal vga_avalon_vga_sink_ready_from_sa : OUT STD_LOGIC;
                 signal vga_avalon_vga_sink_reset : OUT STD_LOGIC;
                 signal vga_avalon_vga_sink_startofpacket : OUT STD_LOGIC;
                 signal vga_avalon_vga_sink_valid : OUT STD_LOGIC
              );
end entity vga_avalon_vga_sink_arbitrator;


architecture europa of vga_avalon_vga_sink_arbitrator is

begin

  --mux vga_avalon_vga_sink_data, which is an e_mux
  vga_avalon_vga_sink_data <= alpha_blending_avalon_blended_source_data;
  --mux vga_avalon_vga_sink_empty, which is an e_mux
  vga_avalon_vga_sink_empty <= alpha_blending_avalon_blended_source_empty;
  --mux vga_avalon_vga_sink_endofpacket, which is an e_mux
  vga_avalon_vga_sink_endofpacket <= alpha_blending_avalon_blended_source_endofpacket;
  --assign vga_avalon_vga_sink_ready_from_sa = vga_avalon_vga_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  vga_avalon_vga_sink_ready_from_sa <= vga_avalon_vga_sink_ready;
  --mux vga_avalon_vga_sink_startofpacket, which is an e_mux
  vga_avalon_vga_sink_startofpacket <= alpha_blending_avalon_blended_source_startofpacket;
  --mux vga_avalon_vga_sink_valid, which is an e_mux
  vga_avalon_vga_sink_valid <= alpha_blending_avalon_blended_source_valid;
  --~vga_avalon_vga_sink_reset assignment, which is an e_assign
  vga_avalon_vga_sink_reset <= NOT reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGAProc_reset_clk_0_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity VGAProc_reset_clk_0_domain_synch_module;


architecture europa of VGAProc_reset_clk_0_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity VGAProc is 
        port (
              -- 1) global signals:
                 signal clk_0 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0
                 signal FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;
                 signal FL_DQ_to_and_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;
                 signal FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;
                 signal FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;

              -- the_analyzer_input_left
                 signal x_in_to_the_analyzer_input_left : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal y_in_to_the_analyzer_input_left : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

              -- the_analyzer_input_right
                 signal x_in_to_the_analyzer_input_right : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal y_in_to_the_analyzer_input_right : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

              -- the_audio_and_video_config_0
                 signal I2C_SCLK_from_the_audio_and_video_config_0 : OUT STD_LOGIC;
                 signal I2C_SDAT_to_and_from_the_audio_and_video_config_0 : INOUT STD_LOGIC;

              -- the_membuffer_0
                 signal delay_time_to_the_membuffer_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sample_clk_to_the_membuffer_0 : IN STD_LOGIC;
                 signal sample_left_in_to_the_membuffer_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sample_left_out_from_the_membuffer_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sample_right_in_to_the_membuffer_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sample_right_out_from_the_membuffer_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_bitcrusher_bypass
                 signal out_port_from_the_pio_bitcrusher_bypass : OUT STD_LOGIC;

              -- the_pio_bitcrusher_crush
                 signal out_port_from_the_pio_bitcrusher_crush : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_pio_bitcrusher_downsample
                 signal out_port_from_the_pio_bitcrusher_downsample : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_pio_bitcrusher_drywet
                 signal out_port_from_the_pio_bitcrusher_drywet : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_bitcrusher_flavor
                 signal out_port_from_the_pio_bitcrusher_flavor : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_pio_bitcrusher_tone
                 signal out_port_from_the_pio_bitcrusher_tone : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_compressor_bypass
                 signal out_port_from_the_pio_compressor_bypass : OUT STD_LOGIC;

              -- the_pio_compressor_gain
                 signal out_port_from_the_pio_compressor_gain : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_pio_compressor_treshold
                 signal out_port_from_the_pio_compressor_treshold : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_delay_bypass
                 signal out_port_from_the_pio_delay_bypass : OUT STD_LOGIC;

              -- the_pio_delay_decay
                 signal out_port_from_the_pio_delay_decay : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_pio_delay_length
                 signal out_port_from_the_pio_delay_length : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_master_volume
                 signal out_port_from_the_pio_master_volume : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_octaver_bypass
                 signal out_port_from_the_pio_octaver_bypass : OUT STD_LOGIC;

              -- the_pio_octaver_dry_wet
                 signal out_port_from_the_pio_octaver_dry_wet : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_output_power_left
                 signal in_port_to_the_pio_output_power_left : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_output_power_right
                 signal in_port_to_the_pio_output_power_right : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_overdrive_asymmetric
                 signal out_port_from_the_pio_overdrive_asymmetric : OUT STD_LOGIC;

              -- the_pio_overdrive_bypass
                 signal out_port_from_the_pio_overdrive_bypass : OUT STD_LOGIC;

              -- the_pio_overdrive_gain
                 signal out_port_from_the_pio_overdrive_gain : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_overdrive_tone
                 signal out_port_from_the_pio_overdrive_tone : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_overdrive_volume
                 signal out_port_from_the_pio_overdrive_volume : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_tremolo_stereo_bypass
                 signal out_port_from_the_pio_tremolo_stereo_bypass : OUT STD_LOGIC;

              -- the_pio_tremolo_stereo_depth
                 signal out_port_from_the_pio_tremolo_stereo_depth : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_pio_tremolo_stereo_mode
                 signal out_port_from_the_pio_tremolo_stereo_mode : OUT STD_LOGIC;

              -- the_pio_tremolo_stereo_sweep_a
                 signal out_port_from_the_pio_tremolo_stereo_sweep_a : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_pio_tremolo_stereo_sweep_b
                 signal out_port_from_the_pio_tremolo_stereo_sweep_b : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_ps2
                 signal PS2_CLK_to_and_from_the_ps2 : INOUT STD_LOGIC;
                 signal PS2_DAT_to_and_from_the_ps2 : INOUT STD_LOGIC;

              -- the_sdram
                 signal zs_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal zs_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_cas_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cke_from_the_sdram : OUT STD_LOGIC;
                 signal zs_cs_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal zs_dqm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_ras_n_from_the_sdram : OUT STD_LOGIC;
                 signal zs_we_n_from_the_sdram : OUT STD_LOGIC;

              -- the_sram
                 signal SRAM_ADDR_from_the_sram : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal SRAM_CE_N_from_the_sram : OUT STD_LOGIC;
                 signal SRAM_DQ_to_and_from_the_sram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal SRAM_LB_N_from_the_sram : OUT STD_LOGIC;
                 signal SRAM_OE_N_from_the_sram : OUT STD_LOGIC;
                 signal SRAM_UB_N_from_the_sram : OUT STD_LOGIC;
                 signal SRAM_WE_N_from_the_sram : OUT STD_LOGIC;

              -- the_vga
                 signal VGA_BLANK_from_the_vga : OUT STD_LOGIC;
                 signal VGA_B_from_the_vga : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal VGA_G_from_the_vga : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal VGA_HS_from_the_vga : OUT STD_LOGIC;
                 signal VGA_R_from_the_vga : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal VGA_SYNC_from_the_vga : OUT STD_LOGIC;
                 signal VGA_VS_from_the_vga : OUT STD_LOGIC
              );
end entity VGAProc;


architecture europa of VGAProc is
component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arbitrator is 
           port (
                 -- inputs:
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                    signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : OUT STD_LOGIC;
                    signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer : OUT STD_LOGIC
                 );
end component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arbitrator;

component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arbitrator is 
           port (
                 -- inputs:
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write : OUT STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                    signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : OUT STD_LOGIC;
                    signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer : OUT STD_LOGIC
                 );
end component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arbitrator;

component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 is 
           port (
                 -- inputs:
                    signal i_avalon_address : IN STD_LOGIC_VECTOR (19 DOWNTO 0);
                    signal i_avalon_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal i_avalon_chip_select : IN STD_LOGIC;
                    signal i_avalon_erase_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal i_avalon_erase_chip_select : IN STD_LOGIC;
                    signal i_avalon_erase_read : IN STD_LOGIC;
                    signal i_avalon_erase_write : IN STD_LOGIC;
                    signal i_avalon_erase_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_avalon_read : IN STD_LOGIC;
                    signal i_avalon_write : IN STD_LOGIC;
                    signal i_avalon_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_clock : IN STD_LOGIC;
                    signal i_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal FL_ADDR : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal FL_CE_N : OUT STD_LOGIC;
                    signal FL_DQ : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal FL_OE_N : OUT STD_LOGIC;
                    signal FL_RST_N : OUT STD_LOGIC;
                    signal FL_WE_N : OUT STD_LOGIC;
                    signal o_avalon_erase_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal o_avalon_erase_waitrequest : OUT STD_LOGIC;
                    signal o_avalon_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal o_avalon_waitrequest : OUT STD_LOGIC
                 );
end component Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0;

component alpha_blending_avalon_background_sink_arbitrator is 
           port (
                 -- inputs:
                    signal alpha_blending_avalon_background_sink_ready : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_source_endofpacket : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_source_startofpacket : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_source_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal alpha_blending_avalon_background_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal alpha_blending_avalon_background_sink_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal alpha_blending_avalon_background_sink_endofpacket : OUT STD_LOGIC;
                    signal alpha_blending_avalon_background_sink_ready_from_sa : OUT STD_LOGIC;
                    signal alpha_blending_avalon_background_sink_startofpacket : OUT STD_LOGIC;
                    signal alpha_blending_avalon_background_sink_valid : OUT STD_LOGIC
                 );
end component alpha_blending_avalon_background_sink_arbitrator;

component alpha_blending_avalon_foreground_sink_arbitrator is 
           port (
                 -- inputs:
                    signal alpha_blending_avalon_foreground_sink_ready : IN STD_LOGIC;
                    signal character_buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal character_buffer_avalon_char_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal character_buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                    signal character_buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                    signal character_buffer_avalon_char_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal alpha_blending_avalon_foreground_sink_data : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal alpha_blending_avalon_foreground_sink_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal alpha_blending_avalon_foreground_sink_endofpacket : OUT STD_LOGIC;
                    signal alpha_blending_avalon_foreground_sink_ready_from_sa : OUT STD_LOGIC;
                    signal alpha_blending_avalon_foreground_sink_reset : OUT STD_LOGIC;
                    signal alpha_blending_avalon_foreground_sink_startofpacket : OUT STD_LOGIC;
                    signal alpha_blending_avalon_foreground_sink_valid : OUT STD_LOGIC
                 );
end component alpha_blending_avalon_foreground_sink_arbitrator;

component alpha_blending_avalon_blended_source_arbitrator is 
           port (
                 -- inputs:
                    signal alpha_blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal alpha_blending_avalon_blended_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal alpha_blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                    signal alpha_blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                    signal alpha_blending_avalon_blended_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal vga_avalon_vga_sink_ready_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal alpha_blending_avalon_blended_source_ready : OUT STD_LOGIC
                 );
end component alpha_blending_avalon_blended_source_arbitrator;

component alpha_blending is 
           port (
                 -- inputs:
                    signal background_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal background_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal background_endofpacket : IN STD_LOGIC;
                    signal background_startofpacket : IN STD_LOGIC;
                    signal background_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal foreground_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal foreground_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal foreground_endofpacket : IN STD_LOGIC;
                    signal foreground_startofpacket : IN STD_LOGIC;
                    signal foreground_valid : IN STD_LOGIC;
                    signal output_ready : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;

                 -- outputs:
                    signal background_ready : OUT STD_LOGIC;
                    signal foreground_ready : OUT STD_LOGIC;
                    signal output_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal output_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal output_endofpacket : OUT STD_LOGIC;
                    signal output_startofpacket : OUT STD_LOGIC;
                    signal output_valid : OUT STD_LOGIC
                 );
end component alpha_blending;

component analyzer_input_left_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal analyzer_input_left_avalon_slave_readdata : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal analyzer_input_left_avalon_slave_read : OUT STD_LOGIC;
                    signal analyzer_input_left_avalon_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
                    signal analyzer_input_left_avalon_slave_reset_n : OUT STD_LOGIC;
                    signal cpu_data_master_granted_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_analyzer_input_left_avalon_slave : OUT STD_LOGIC;
                    signal d1_analyzer_input_left_avalon_slave_end_xfer : OUT STD_LOGIC
                 );
end component analyzer_input_left_avalon_slave_arbitrator;

component analyzer_input_left is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal x_in : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal y_in : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (127 DOWNTO 0)
                 );
end component analyzer_input_left;

component analyzer_input_right_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal analyzer_input_right_avalon_slave_readdata : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal analyzer_input_right_avalon_slave_read : OUT STD_LOGIC;
                    signal analyzer_input_right_avalon_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
                    signal analyzer_input_right_avalon_slave_reset_n : OUT STD_LOGIC;
                    signal cpu_data_master_granted_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_analyzer_input_right_avalon_slave : OUT STD_LOGIC;
                    signal d1_analyzer_input_right_avalon_slave_end_xfer : OUT STD_LOGIC
                 );
end component analyzer_input_right_avalon_slave_arbitrator;

component analyzer_input_right is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal x_in : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal y_in : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (127 DOWNTO 0)
                 );
end component analyzer_input_right;

component audio_and_video_config_0_avalon_on_board_config_slave_arbitrator is 
           port (
                 -- inputs:
                    signal audio_and_video_config_0_avalon_on_board_config_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal audio_and_video_config_0_avalon_on_board_config_slave_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal audio_and_video_config_0_avalon_on_board_config_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal audio_and_video_config_0_avalon_on_board_config_slave_chipselect : OUT STD_LOGIC;
                    signal audio_and_video_config_0_avalon_on_board_config_slave_read : OUT STD_LOGIC;
                    signal audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal audio_and_video_config_0_avalon_on_board_config_slave_reset : OUT STD_LOGIC;
                    signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal audio_and_video_config_0_avalon_on_board_config_slave_write : OUT STD_LOGIC;
                    signal audio_and_video_config_0_avalon_on_board_config_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC;
                    signal d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : OUT STD_LOGIC
                 );
end component audio_and_video_config_0_avalon_on_board_config_slave_arbitrator;

component audio_and_video_config_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal ob_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal ob_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ob_chipselect : IN STD_LOGIC;
                    signal ob_read : IN STD_LOGIC;
                    signal ob_write : IN STD_LOGIC;
                    signal ob_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset : IN STD_LOGIC;

                 -- outputs:
                    signal I2C_SCLK : OUT STD_LOGIC;
                    signal I2C_SDAT : INOUT STD_LOGIC;
                    signal ob_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ob_waitrequest : OUT STD_LOGIC
                 );
end component audio_and_video_config_0;

component character_buffer_avalon_char_buffer_slave_arbitrator is 
           port (
                 -- inputs:
                    signal character_buffer_avalon_char_buffer_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal character_buffer_avalon_char_buffer_slave_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal character_buffer_avalon_char_buffer_slave_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal character_buffer_avalon_char_buffer_slave_chipselect : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_buffer_slave_read : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_buffer_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal character_buffer_avalon_char_buffer_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_buffer_slave_write : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_buffer_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal cpu_data_master_granted_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC;
                    signal d1_character_buffer_avalon_char_buffer_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : OUT STD_LOGIC
                 );
end component character_buffer_avalon_char_buffer_slave_arbitrator;

component character_buffer_avalon_char_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal character_buffer_avalon_char_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal character_buffer_avalon_char_control_slave_address : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_control_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal character_buffer_avalon_char_control_slave_chipselect : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_control_slave_read : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal character_buffer_avalon_char_control_slave_reset : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_control_slave_write : OUT STD_LOGIC;
                    signal character_buffer_avalon_char_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_granted_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_character_buffer_avalon_char_control_slave : OUT STD_LOGIC;
                    signal d1_character_buffer_avalon_char_control_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : OUT STD_LOGIC
                 );
end component character_buffer_avalon_char_control_slave_arbitrator;

component character_buffer_avalon_char_source_arbitrator is 
           port (
                 -- inputs:
                    signal alpha_blending_avalon_foreground_sink_ready_from_sa : IN STD_LOGIC;
                    signal character_buffer_avalon_char_source_data : IN STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal character_buffer_avalon_char_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal character_buffer_avalon_char_source_endofpacket : IN STD_LOGIC;
                    signal character_buffer_avalon_char_source_startofpacket : IN STD_LOGIC;
                    signal character_buffer_avalon_char_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal character_buffer_avalon_char_source_ready : OUT STD_LOGIC
                 );
end component character_buffer_avalon_char_source_arbitrator;

component character_buffer is 
           port (
                 -- inputs:
                    signal buf_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal buf_chipselect : IN STD_LOGIC;
                    signal buf_read : IN STD_LOGIC;
                    signal buf_write : IN STD_LOGIC;
                    signal buf_writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal ctrl_address : IN STD_LOGIC;
                    signal ctrl_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ctrl_chipselect : IN STD_LOGIC;
                    signal ctrl_read : IN STD_LOGIC;
                    signal ctrl_write : IN STD_LOGIC;
                    signal ctrl_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset : IN STD_LOGIC;
                    signal stream_ready : IN STD_LOGIC;

                 -- outputs:
                    signal buf_readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal buf_waitrequest : OUT STD_LOGIC;
                    signal ctrl_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal stream_data : OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
                    signal stream_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal stream_endofpacket : OUT STD_LOGIC;
                    signal stream_startofpacket : OUT STD_LOGIC;
                    signal stream_valid : OUT STD_LOGIC
                 );
end component character_buffer;

component cpu_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_data_master_requests_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_instruction_master_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_write : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC
                 );
end component cpu_jtag_debug_module_arbitrator;

component cpu_custom_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_custom_instruction_master_multi_start : IN STD_LOGIC;
                    signal cpu_fpoint_s1_done_from_sa : IN STD_LOGIC;
                    signal cpu_fpoint_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_custom_instruction_master_multi_done : OUT STD_LOGIC;
                    signal cpu_custom_instruction_master_multi_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_custom_instruction_master_reset_n : OUT STD_LOGIC;
                    signal cpu_custom_instruction_master_start_cpu_fpoint_s1 : OUT STD_LOGIC;
                    signal cpu_fpoint_s1_select : OUT STD_LOGIC
                 );
end component cpu_custom_instruction_master_arbitrator;

component cpu_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa : IN STD_LOGIC;
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa : IN STD_LOGIC;
                    signal analyzer_input_left_avalon_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                    signal analyzer_input_right_avalon_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
                    signal audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal character_buffer_avalon_char_buffer_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal character_buffer_avalon_char_buffer_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal character_buffer_avalon_char_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_byteenable_sdram_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_byteenable_sram_avalon_sram_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                    signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                    signal cpu_data_master_granted_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_data_master_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_compressor_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_compressor_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_compressor_treshold_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_delay_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_delay_decay_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_delay_length_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_master_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_octaver_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_output_power_left_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_output_power_right_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_overdrive_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_overdrive_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_overdrive_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_ps2_avalon_ps2_slave : IN STD_LOGIC;
                    signal cpu_data_master_granted_sdram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_compressor_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_compressor_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_compressor_treshold_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_delay_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_delay_decay_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_delay_length_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_master_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_octaver_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_output_power_left_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_output_power_right_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_ps2_avalon_ps2_slave : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_compressor_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_compressor_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_compressor_treshold_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_delay_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_delay_decay_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_delay_length_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_master_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_octaver_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_output_power_left_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_output_power_right_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : IN STD_LOGIC;
                    signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : IN STD_LOGIC;
                    signal cpu_data_master_requests_analyzer_input_left_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_analyzer_input_right_avalon_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_data_master_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_crush_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_downsample_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_drywet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_flavor_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_compressor_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_compressor_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_compressor_treshold_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_delay_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_delay_decay_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_delay_length_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_master_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_octaver_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_octaver_dry_wet_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_output_power_left_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_output_power_right_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_asymmetric_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_gain_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_tone_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_volume_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_depth_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_mode_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_ps2_avalon_ps2_slave : IN STD_LOGIC;
                    signal cpu_data_master_requests_sdram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer : IN STD_LOGIC;
                    signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer : IN STD_LOGIC;
                    signal d1_analyzer_input_left_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal d1_analyzer_input_right_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer : IN STD_LOGIC;
                    signal d1_character_buffer_avalon_char_buffer_slave_end_xfer : IN STD_LOGIC;
                    signal d1_character_buffer_avalon_char_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal d1_pio_bitcrusher_bypass_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_bitcrusher_crush_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_bitcrusher_downsample_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_bitcrusher_drywet_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_bitcrusher_flavor_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_bitcrusher_tone_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_compressor_bypass_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_compressor_gain_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_compressor_treshold_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_delay_bypass_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_delay_decay_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_delay_length_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_master_volume_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_octaver_bypass_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_octaver_dry_wet_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_output_power_left_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_output_power_right_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_overdrive_asymmetric_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_overdrive_bypass_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_overdrive_gain_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_overdrive_tone_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_overdrive_volume_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_tremolo_stereo_bypass_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_tremolo_stereo_depth_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_tremolo_stereo_mode_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_tremolo_stereo_sweep_a_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pio_tremolo_stereo_sweep_b_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer : IN STD_LOGIC;
                    signal d1_ps2_avalon_ps2_slave_end_xfer : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sram_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal pio_bitcrusher_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_bitcrusher_crush_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pio_bitcrusher_downsample_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pio_bitcrusher_drywet_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_bitcrusher_flavor_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pio_bitcrusher_tone_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_compressor_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_compressor_gain_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pio_compressor_treshold_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_delay_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_delay_decay_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pio_delay_length_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_master_volume_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_octaver_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_octaver_dry_wet_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_output_power_left_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_output_power_right_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_overdrive_asymmetric_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_overdrive_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_overdrive_gain_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_overdrive_tone_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_overdrive_volume_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_tremolo_stereo_bypass_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_tremolo_stereo_depth_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_tremolo_stereo_mode_s1_readdata_from_sa : IN STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_a_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pio_tremolo_stereo_sweep_b_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ps2_avalon_ps2_slave_irq_from_sa : IN STD_LOGIC;
                    signal ps2_avalon_ps2_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ps2_avalon_ps2_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave : IN STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave : IN STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave : IN STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : IN STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : IN STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal sram_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_data_master_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_no_byte_enables_and_last_term : OUT STD_LOGIC;
                    signal cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_data_master_arbitrator;

component cpu_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_instruction_master_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_instruction_master_granted_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_sram_avalon_sram_slave : IN STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_sram_avalon_sram_slave_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sram_avalon_sram_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal cpu_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_instruction_master_arbitrator;

component cpu is 
           port (
                 -- inputs:
                    signal A_ci_multi_done : IN STD_LOGIC;
                    signal A_ci_multi_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal A_ci_multi_a : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal A_ci_multi_b : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal A_ci_multi_c : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal A_ci_multi_clk_en : OUT STD_LOGIC;
                    signal A_ci_multi_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal A_ci_multi_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal A_ci_multi_estatus : OUT STD_LOGIC;
                    signal A_ci_multi_ipending : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal A_ci_multi_n : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal A_ci_multi_readra : OUT STD_LOGIC;
                    signal A_ci_multi_readrb : OUT STD_LOGIC;
                    signal A_ci_multi_start : OUT STD_LOGIC;
                    signal A_ci_multi_status : OUT STD_LOGIC;
                    signal A_ci_multi_writerc : OUT STD_LOGIC;
                    signal d_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component cpu;

component cpu_fpoint_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_custom_instruction_master_multi_clk_en : IN STD_LOGIC;
                    signal cpu_custom_instruction_master_multi_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_custom_instruction_master_multi_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_custom_instruction_master_multi_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal cpu_custom_instruction_master_start_cpu_fpoint_s1 : IN STD_LOGIC;
                    signal cpu_fpoint_s1_done : IN STD_LOGIC;
                    signal cpu_fpoint_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_fpoint_s1_select : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_fpoint_s1_clk_en : OUT STD_LOGIC;
                    signal cpu_fpoint_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_fpoint_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_fpoint_s1_done_from_sa : OUT STD_LOGIC;
                    signal cpu_fpoint_s1_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_fpoint_s1_reset : OUT STD_LOGIC;
                    signal cpu_fpoint_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_fpoint_s1_start : OUT STD_LOGIC
                 );
end component cpu_fpoint_s1_arbitrator;

component cpu_fpoint is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clk_en : IN STD_LOGIC;
                    signal dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reset : IN STD_LOGIC;
                    signal start : IN STD_LOGIC;

                 -- outputs:
                    signal done : OUT STD_LOGIC;
                    signal result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component cpu_fpoint;

component jtag_uart_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component jtag_uart_avalon_jtag_slave_arbitrator;

component jtag_uart is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart;

component membuffer_0_avalon_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal membuffer_0_avalon_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal membuffer_0_avalon_master_read : IN STD_LOGIC;
                    signal membuffer_0_avalon_master_write : IN STD_LOGIC;
                    signal membuffer_0_avalon_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal membuffer_0_byteenable_sdram_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal membuffer_0_granted_sdram_s1 : IN STD_LOGIC;
                    signal membuffer_0_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal membuffer_0_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal membuffer_0_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal membuffer_0_requests_sdram_s1 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal membuffer_0_avalon_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal membuffer_0_avalon_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal membuffer_0_avalon_master_reset_n : OUT STD_LOGIC;
                    signal membuffer_0_avalon_master_waitrequest : OUT STD_LOGIC;
                    signal membuffer_0_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal membuffer_0_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component membuffer_0_avalon_master_arbitrator;

component membuffer_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal delay_time : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset : IN STD_LOGIC;
                    signal sample_clk : IN STD_LOGIC;
                    signal sample_left_in : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sample_right_in : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal read : OUT STD_LOGIC;
                    signal sample_left_out : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sample_right_out : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal write : OUT STD_LOGIC;
                    signal writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component membuffer_0;

component pio_bitcrusher_bypass_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_bitcrusher_bypass_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_bypass_s1 : OUT STD_LOGIC;
                    signal d1_pio_bitcrusher_bypass_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_bitcrusher_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_bitcrusher_bypass_s1_chipselect : OUT STD_LOGIC;
                    signal pio_bitcrusher_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_bitcrusher_bypass_s1_reset_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_bypass_s1_write_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_bypass_s1_writedata : OUT STD_LOGIC
                 );
end component pio_bitcrusher_bypass_s1_arbitrator;

component pio_bitcrusher_bypass is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_bitcrusher_bypass;

component pio_bitcrusher_crush_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_bitcrusher_crush_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_crush_s1 : OUT STD_LOGIC;
                    signal d1_pio_bitcrusher_crush_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_bitcrusher_crush_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_bitcrusher_crush_s1_chipselect : OUT STD_LOGIC;
                    signal pio_bitcrusher_crush_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pio_bitcrusher_crush_s1_reset_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_crush_s1_write_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_crush_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_bitcrusher_crush_s1_arbitrator;

component pio_bitcrusher_crush is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_bitcrusher_crush;

component pio_bitcrusher_downsample_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_bitcrusher_downsample_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_downsample_s1 : OUT STD_LOGIC;
                    signal d1_pio_bitcrusher_downsample_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_bitcrusher_downsample_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_bitcrusher_downsample_s1_chipselect : OUT STD_LOGIC;
                    signal pio_bitcrusher_downsample_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pio_bitcrusher_downsample_s1_reset_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_downsample_s1_write_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_downsample_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component pio_bitcrusher_downsample_s1_arbitrator;

component pio_bitcrusher_downsample is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component pio_bitcrusher_downsample;

component pio_bitcrusher_drywet_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_bitcrusher_drywet_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_drywet_s1 : OUT STD_LOGIC;
                    signal d1_pio_bitcrusher_drywet_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_bitcrusher_drywet_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_bitcrusher_drywet_s1_chipselect : OUT STD_LOGIC;
                    signal pio_bitcrusher_drywet_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_bitcrusher_drywet_s1_reset_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_drywet_s1_write_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_drywet_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_bitcrusher_drywet_s1_arbitrator;

component pio_bitcrusher_drywet is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_bitcrusher_drywet;

component pio_bitcrusher_flavor_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_bitcrusher_flavor_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_flavor_s1 : OUT STD_LOGIC;
                    signal d1_pio_bitcrusher_flavor_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_bitcrusher_flavor_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_bitcrusher_flavor_s1_chipselect : OUT STD_LOGIC;
                    signal pio_bitcrusher_flavor_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pio_bitcrusher_flavor_s1_reset_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_flavor_s1_write_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_flavor_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_bitcrusher_flavor_s1_arbitrator;

component pio_bitcrusher_flavor is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_bitcrusher_flavor;

component pio_bitcrusher_tone_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_bitcrusher_tone_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_bitcrusher_tone_s1 : OUT STD_LOGIC;
                    signal d1_pio_bitcrusher_tone_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_bitcrusher_tone_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_bitcrusher_tone_s1_chipselect : OUT STD_LOGIC;
                    signal pio_bitcrusher_tone_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_bitcrusher_tone_s1_reset_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_tone_s1_write_n : OUT STD_LOGIC;
                    signal pio_bitcrusher_tone_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_bitcrusher_tone_s1_arbitrator;

component pio_bitcrusher_tone is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_bitcrusher_tone;

component pio_compressor_bypass_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_compressor_bypass_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_compressor_bypass_s1 : OUT STD_LOGIC;
                    signal d1_pio_compressor_bypass_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_compressor_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_compressor_bypass_s1_chipselect : OUT STD_LOGIC;
                    signal pio_compressor_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_compressor_bypass_s1_reset_n : OUT STD_LOGIC;
                    signal pio_compressor_bypass_s1_write_n : OUT STD_LOGIC;
                    signal pio_compressor_bypass_s1_writedata : OUT STD_LOGIC
                 );
end component pio_compressor_bypass_s1_arbitrator;

component pio_compressor_bypass is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_compressor_bypass;

component pio_compressor_gain_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_compressor_gain_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_compressor_gain_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_compressor_gain_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_compressor_gain_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_compressor_gain_s1 : OUT STD_LOGIC;
                    signal d1_pio_compressor_gain_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_compressor_gain_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_compressor_gain_s1_chipselect : OUT STD_LOGIC;
                    signal pio_compressor_gain_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pio_compressor_gain_s1_reset_n : OUT STD_LOGIC;
                    signal pio_compressor_gain_s1_write_n : OUT STD_LOGIC;
                    signal pio_compressor_gain_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component pio_compressor_gain_s1_arbitrator;

component pio_compressor_gain is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component pio_compressor_gain;

component pio_compressor_treshold_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_compressor_treshold_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_compressor_treshold_s1 : OUT STD_LOGIC;
                    signal d1_pio_compressor_treshold_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_compressor_treshold_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_compressor_treshold_s1_chipselect : OUT STD_LOGIC;
                    signal pio_compressor_treshold_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_compressor_treshold_s1_reset_n : OUT STD_LOGIC;
                    signal pio_compressor_treshold_s1_write_n : OUT STD_LOGIC;
                    signal pio_compressor_treshold_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_compressor_treshold_s1_arbitrator;

component pio_compressor_treshold is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_compressor_treshold;

component pio_delay_bypass_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_delay_bypass_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_delay_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_delay_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_delay_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_delay_bypass_s1 : OUT STD_LOGIC;
                    signal d1_pio_delay_bypass_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_delay_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_delay_bypass_s1_chipselect : OUT STD_LOGIC;
                    signal pio_delay_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_delay_bypass_s1_reset_n : OUT STD_LOGIC;
                    signal pio_delay_bypass_s1_write_n : OUT STD_LOGIC;
                    signal pio_delay_bypass_s1_writedata : OUT STD_LOGIC
                 );
end component pio_delay_bypass_s1_arbitrator;

component pio_delay_bypass is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_delay_bypass;

component pio_delay_decay_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_delay_decay_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_delay_decay_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_delay_decay_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_delay_decay_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_delay_decay_s1 : OUT STD_LOGIC;
                    signal d1_pio_delay_decay_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_delay_decay_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_delay_decay_s1_chipselect : OUT STD_LOGIC;
                    signal pio_delay_decay_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pio_delay_decay_s1_reset_n : OUT STD_LOGIC;
                    signal pio_delay_decay_s1_write_n : OUT STD_LOGIC;
                    signal pio_delay_decay_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component pio_delay_decay_s1_arbitrator;

component pio_delay_decay is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component pio_delay_decay;

component pio_delay_length_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_delay_length_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_delay_length_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_delay_length_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_delay_length_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_delay_length_s1 : OUT STD_LOGIC;
                    signal d1_pio_delay_length_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_delay_length_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_delay_length_s1_chipselect : OUT STD_LOGIC;
                    signal pio_delay_length_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_delay_length_s1_reset_n : OUT STD_LOGIC;
                    signal pio_delay_length_s1_write_n : OUT STD_LOGIC;
                    signal pio_delay_length_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_delay_length_s1_arbitrator;

component pio_delay_length is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_delay_length;

component pio_master_volume_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_master_volume_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_master_volume_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_master_volume_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_master_volume_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_master_volume_s1 : OUT STD_LOGIC;
                    signal d1_pio_master_volume_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_master_volume_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_master_volume_s1_chipselect : OUT STD_LOGIC;
                    signal pio_master_volume_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_master_volume_s1_reset_n : OUT STD_LOGIC;
                    signal pio_master_volume_s1_write_n : OUT STD_LOGIC;
                    signal pio_master_volume_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_master_volume_s1_arbitrator;

component pio_master_volume is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_master_volume;

component pio_octaver_bypass_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_octaver_bypass_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_octaver_bypass_s1 : OUT STD_LOGIC;
                    signal d1_pio_octaver_bypass_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_octaver_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_octaver_bypass_s1_chipselect : OUT STD_LOGIC;
                    signal pio_octaver_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_octaver_bypass_s1_reset_n : OUT STD_LOGIC;
                    signal pio_octaver_bypass_s1_write_n : OUT STD_LOGIC;
                    signal pio_octaver_bypass_s1_writedata : OUT STD_LOGIC
                 );
end component pio_octaver_bypass_s1_arbitrator;

component pio_octaver_bypass is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_octaver_bypass;

component pio_octaver_dry_wet_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_octaver_dry_wet_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_octaver_dry_wet_s1 : OUT STD_LOGIC;
                    signal d1_pio_octaver_dry_wet_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_octaver_dry_wet_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_octaver_dry_wet_s1_chipselect : OUT STD_LOGIC;
                    signal pio_octaver_dry_wet_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_octaver_dry_wet_s1_reset_n : OUT STD_LOGIC;
                    signal pio_octaver_dry_wet_s1_write_n : OUT STD_LOGIC;
                    signal pio_octaver_dry_wet_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_octaver_dry_wet_s1_arbitrator;

component pio_octaver_dry_wet is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_octaver_dry_wet;

component pio_output_power_left_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal pio_output_power_left_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_output_power_left_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_output_power_left_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_output_power_left_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_output_power_left_s1 : OUT STD_LOGIC;
                    signal d1_pio_output_power_left_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_output_power_left_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_output_power_left_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_output_power_left_s1_reset_n : OUT STD_LOGIC
                 );
end component pio_output_power_left_s1_arbitrator;

component pio_output_power_left is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_output_power_left;

component pio_output_power_right_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal pio_output_power_right_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_output_power_right_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_output_power_right_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_output_power_right_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_output_power_right_s1 : OUT STD_LOGIC;
                    signal d1_pio_output_power_right_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_output_power_right_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_output_power_right_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_output_power_right_s1_reset_n : OUT STD_LOGIC
                 );
end component pio_output_power_right_s1_arbitrator;

component pio_output_power_right is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_output_power_right;

component pio_overdrive_asymmetric_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_overdrive_asymmetric_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_asymmetric_s1 : OUT STD_LOGIC;
                    signal d1_pio_overdrive_asymmetric_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_overdrive_asymmetric_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_overdrive_asymmetric_s1_chipselect : OUT STD_LOGIC;
                    signal pio_overdrive_asymmetric_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_overdrive_asymmetric_s1_reset_n : OUT STD_LOGIC;
                    signal pio_overdrive_asymmetric_s1_write_n : OUT STD_LOGIC;
                    signal pio_overdrive_asymmetric_s1_writedata : OUT STD_LOGIC
                 );
end component pio_overdrive_asymmetric_s1_arbitrator;

component pio_overdrive_asymmetric is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_overdrive_asymmetric;

component pio_overdrive_bypass_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_overdrive_bypass_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_bypass_s1 : OUT STD_LOGIC;
                    signal d1_pio_overdrive_bypass_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_overdrive_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_overdrive_bypass_s1_chipselect : OUT STD_LOGIC;
                    signal pio_overdrive_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_overdrive_bypass_s1_reset_n : OUT STD_LOGIC;
                    signal pio_overdrive_bypass_s1_write_n : OUT STD_LOGIC;
                    signal pio_overdrive_bypass_s1_writedata : OUT STD_LOGIC
                 );
end component pio_overdrive_bypass_s1_arbitrator;

component pio_overdrive_bypass is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_overdrive_bypass;

component pio_overdrive_gain_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_overdrive_gain_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_gain_s1 : OUT STD_LOGIC;
                    signal d1_pio_overdrive_gain_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_overdrive_gain_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_overdrive_gain_s1_chipselect : OUT STD_LOGIC;
                    signal pio_overdrive_gain_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_overdrive_gain_s1_reset_n : OUT STD_LOGIC;
                    signal pio_overdrive_gain_s1_write_n : OUT STD_LOGIC;
                    signal pio_overdrive_gain_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_overdrive_gain_s1_arbitrator;

component pio_overdrive_gain is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_overdrive_gain;

component pio_overdrive_tone_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_overdrive_tone_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_tone_s1 : OUT STD_LOGIC;
                    signal d1_pio_overdrive_tone_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_overdrive_tone_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_overdrive_tone_s1_chipselect : OUT STD_LOGIC;
                    signal pio_overdrive_tone_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_overdrive_tone_s1_reset_n : OUT STD_LOGIC;
                    signal pio_overdrive_tone_s1_write_n : OUT STD_LOGIC;
                    signal pio_overdrive_tone_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_overdrive_tone_s1_arbitrator;

component pio_overdrive_tone is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_overdrive_tone;

component pio_overdrive_volume_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_overdrive_volume_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_overdrive_volume_s1 : OUT STD_LOGIC;
                    signal d1_pio_overdrive_volume_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_overdrive_volume_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_overdrive_volume_s1_chipselect : OUT STD_LOGIC;
                    signal pio_overdrive_volume_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_overdrive_volume_s1_reset_n : OUT STD_LOGIC;
                    signal pio_overdrive_volume_s1_write_n : OUT STD_LOGIC;
                    signal pio_overdrive_volume_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_overdrive_volume_s1_arbitrator;

component pio_overdrive_volume is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_overdrive_volume;

component pio_tremolo_stereo_bypass_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_tremolo_stereo_bypass_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 : OUT STD_LOGIC;
                    signal d1_pio_tremolo_stereo_bypass_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_bypass_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_tremolo_stereo_bypass_s1_chipselect : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_bypass_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_bypass_s1_reset_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_bypass_s1_write_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_bypass_s1_writedata : OUT STD_LOGIC
                 );
end component pio_tremolo_stereo_bypass_s1_arbitrator;

component pio_tremolo_stereo_bypass is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_tremolo_stereo_bypass;

component pio_tremolo_stereo_depth_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_tremolo_stereo_depth_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_depth_s1 : OUT STD_LOGIC;
                    signal d1_pio_tremolo_stereo_depth_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_depth_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_tremolo_stereo_depth_s1_chipselect : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_depth_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pio_tremolo_stereo_depth_s1_reset_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_depth_s1_write_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_depth_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_tremolo_stereo_depth_s1_arbitrator;

component pio_tremolo_stereo_depth is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pio_tremolo_stereo_depth;

component pio_tremolo_stereo_mode_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_tremolo_stereo_mode_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_mode_s1 : OUT STD_LOGIC;
                    signal d1_pio_tremolo_stereo_mode_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_mode_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_tremolo_stereo_mode_s1_chipselect : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_mode_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_mode_s1_reset_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_mode_s1_write_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_mode_s1_writedata : OUT STD_LOGIC
                 );
end component pio_tremolo_stereo_mode_s1_arbitrator;

component pio_tremolo_stereo_mode is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component pio_tremolo_stereo_mode;

component pio_tremolo_stereo_sweep_a_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_tremolo_stereo_sweep_a_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 : OUT STD_LOGIC;
                    signal d1_pio_tremolo_stereo_sweep_a_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_a_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_tremolo_stereo_sweep_a_s1_chipselect : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_a_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pio_tremolo_stereo_sweep_a_s1_reset_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_a_s1_write_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_a_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_tremolo_stereo_sweep_a_s1_arbitrator;

component pio_tremolo_stereo_sweep_a is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_tremolo_stereo_sweep_a;

component pio_tremolo_stereo_sweep_b_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pio_tremolo_stereo_sweep_b_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 : OUT STD_LOGIC;
                    signal d1_pio_tremolo_stereo_sweep_b_s1_end_xfer : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_b_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pio_tremolo_stereo_sweep_b_s1_chipselect : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_b_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pio_tremolo_stereo_sweep_b_s1_reset_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_b_s1_write_n : OUT STD_LOGIC;
                    signal pio_tremolo_stereo_sweep_b_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_tremolo_stereo_sweep_b_s1_arbitrator;

component pio_tremolo_stereo_sweep_b is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component pio_tremolo_stereo_sweep_b;

component pixel_buffer_avalon_pixel_buffer_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC;
                    signal d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_slave_read : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_slave_reset : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_slave_write : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave : OUT STD_LOGIC
                 );
end component pixel_buffer_avalon_pixel_buffer_slave_arbitrator;

component pixel_buffer_avalon_pixel_buffer_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_read : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal pixel_buffer_avalon_pixel_buffer_master_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_master_latency_counter : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_master_readdatavalid : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_waitrequest : OUT STD_LOGIC
                 );
end component pixel_buffer_avalon_pixel_buffer_master_arbitrator;

component pixel_buffer_avalon_pixel_buffer_source_arbitrator is 
           port (
                 -- inputs:
                    signal alpha_blending_avalon_background_sink_ready_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_source_endofpacket : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_source_startofpacket : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_source_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pixel_buffer_avalon_pixel_buffer_source_ready : OUT STD_LOGIC
                 );
end component pixel_buffer_avalon_pixel_buffer_source_arbitrator;

component pixel_buffer is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal stream_ready : IN STD_LOGIC;

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_arbiterlock : OUT STD_LOGIC;
                    signal master_read : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal stream_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal stream_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal stream_endofpacket : OUT STD_LOGIC;
                    signal stream_startofpacket : OUT STD_LOGIC;
                    signal stream_valid : OUT STD_LOGIC
                 );
end component pixel_buffer;

component ps2_avalon_ps2_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ps2_avalon_ps2_slave_irq : IN STD_LOGIC;
                    signal ps2_avalon_ps2_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ps2_avalon_ps2_slave_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_ps2_avalon_ps2_slave : OUT STD_LOGIC;
                    signal d1_ps2_avalon_ps2_slave_end_xfer : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_address : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ps2_avalon_ps2_slave_chipselect : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_irq_from_sa : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_read : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ps2_avalon_ps2_slave_reset : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_write : OUT STD_LOGIC;
                    signal ps2_avalon_ps2_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave : OUT STD_LOGIC
                 );
end component ps2_avalon_ps2_slave_arbitrator;

component ps2 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal PS2_CLK : INOUT STD_LOGIC;
                    signal PS2_DAT : INOUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component ps2;

component sdram_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal membuffer_0_avalon_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal membuffer_0_avalon_master_read : IN STD_LOGIC;
                    signal membuffer_0_avalon_master_write : IN STD_LOGIC;
                    signal membuffer_0_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal membuffer_0_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_master_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pixel_buffer_avalon_pixel_buffer_master_arbiterlock : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_latency_counter : IN STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_readdatavalid : IN STD_LOGIC;
                    signal sdram_s1_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_byteenable_sdram_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_granted_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_sdram_s1 : OUT STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                    signal membuffer_0_byteenable_sdram_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal membuffer_0_granted_sdram_s1 : OUT STD_LOGIC;
                    signal membuffer_0_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal membuffer_0_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal membuffer_0_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal membuffer_0_requests_sdram_s1 : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 : OUT STD_LOGIC;
                    signal sdram_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal sdram_s1_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sdram_s1_chipselect : OUT STD_LOGIC;
                    signal sdram_s1_read_n : OUT STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sdram_s1_reset_n : OUT STD_LOGIC;
                    signal sdram_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal sdram_s1_write_n : OUT STD_LOGIC;
                    signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sdram_s1_arbitrator;

component sdram is 
           port (
                 -- inputs:
                    signal az_addr : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal az_be_n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal az_cs : IN STD_LOGIC;
                    signal az_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal az_rd_n : IN STD_LOGIC;
                    signal az_wr_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal za_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal za_valid : OUT STD_LOGIC;
                    signal za_waitrequest : OUT STD_LOGIC;
                    signal zs_addr : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : OUT STD_LOGIC;
                    signal zs_cke : OUT STD_LOGIC;
                    signal zs_cs_n : OUT STD_LOGIC;
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n : OUT STD_LOGIC;
                    signal zs_we_n : OUT STD_LOGIC
                 );
end component sdram;

component sram_avalon_sram_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sram_avalon_sram_slave_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal cpu_data_master_byteenable_sram_avalon_sram_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cpu_data_master_granted_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal cpu_data_master_requests_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal cpu_instruction_master_granted_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal d1_sram_avalon_sram_slave_end_xfer : OUT STD_LOGIC;
                    signal registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave : OUT STD_LOGIC;
                    signal sram_avalon_sram_slave_address : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal sram_avalon_sram_slave_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sram_avalon_sram_slave_read : OUT STD_LOGIC;
                    signal sram_avalon_sram_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sram_avalon_sram_slave_reset : OUT STD_LOGIC;
                    signal sram_avalon_sram_slave_write : OUT STD_LOGIC;
                    signal sram_avalon_sram_slave_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sram_avalon_sram_slave_arbitrator;

component sram is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal SRAM_ADDR : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal SRAM_CE_N : OUT STD_LOGIC;
                    signal SRAM_DQ : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SRAM_LB_N : OUT STD_LOGIC;
                    signal SRAM_OE_N : OUT STD_LOGIC;
                    signal SRAM_UB_N : OUT STD_LOGIC;
                    signal SRAM_WE_N : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sram;

component vga_avalon_vga_sink_arbitrator is 
           port (
                 -- inputs:
                    signal alpha_blending_avalon_blended_source_data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal alpha_blending_avalon_blended_source_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal alpha_blending_avalon_blended_source_endofpacket : IN STD_LOGIC;
                    signal alpha_blending_avalon_blended_source_startofpacket : IN STD_LOGIC;
                    signal alpha_blending_avalon_blended_source_valid : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal vga_avalon_vga_sink_ready : IN STD_LOGIC;

                 -- outputs:
                    signal vga_avalon_vga_sink_data : OUT STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal vga_avalon_vga_sink_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal vga_avalon_vga_sink_endofpacket : OUT STD_LOGIC;
                    signal vga_avalon_vga_sink_ready_from_sa : OUT STD_LOGIC;
                    signal vga_avalon_vga_sink_reset : OUT STD_LOGIC;
                    signal vga_avalon_vga_sink_startofpacket : OUT STD_LOGIC;
                    signal vga_avalon_vga_sink_valid : OUT STD_LOGIC
                 );
end component vga_avalon_vga_sink_arbitrator;

component vga is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (29 DOWNTO 0);
                    signal empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal endofpacket : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal startofpacket : IN STD_LOGIC;
                    signal valid : IN STD_LOGIC;

                 -- outputs:
                    signal VGA_B : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_BLANK : OUT STD_LOGIC;
                    signal VGA_G : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_HS : OUT STD_LOGIC;
                    signal VGA_R : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_SYNC : OUT STD_LOGIC;
                    signal VGA_VS : OUT STD_LOGIC;
                    signal ready : OUT STD_LOGIC
                 );
end component vga;

component VGAProc_reset_clk_0_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component VGAProc_reset_clk_0_domain_synch_module;

                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address :  STD_LOGIC_VECTOR (19 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write :  STD_LOGIC;
                signal Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal alpha_blending_avalon_background_sink_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal alpha_blending_avalon_background_sink_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal alpha_blending_avalon_background_sink_endofpacket :  STD_LOGIC;
                signal alpha_blending_avalon_background_sink_ready :  STD_LOGIC;
                signal alpha_blending_avalon_background_sink_ready_from_sa :  STD_LOGIC;
                signal alpha_blending_avalon_background_sink_startofpacket :  STD_LOGIC;
                signal alpha_blending_avalon_background_sink_valid :  STD_LOGIC;
                signal alpha_blending_avalon_blended_source_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal alpha_blending_avalon_blended_source_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal alpha_blending_avalon_blended_source_endofpacket :  STD_LOGIC;
                signal alpha_blending_avalon_blended_source_ready :  STD_LOGIC;
                signal alpha_blending_avalon_blended_source_startofpacket :  STD_LOGIC;
                signal alpha_blending_avalon_blended_source_valid :  STD_LOGIC;
                signal alpha_blending_avalon_foreground_sink_data :  STD_LOGIC_VECTOR (39 DOWNTO 0);
                signal alpha_blending_avalon_foreground_sink_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal alpha_blending_avalon_foreground_sink_endofpacket :  STD_LOGIC;
                signal alpha_blending_avalon_foreground_sink_ready :  STD_LOGIC;
                signal alpha_blending_avalon_foreground_sink_ready_from_sa :  STD_LOGIC;
                signal alpha_blending_avalon_foreground_sink_reset :  STD_LOGIC;
                signal alpha_blending_avalon_foreground_sink_startofpacket :  STD_LOGIC;
                signal alpha_blending_avalon_foreground_sink_valid :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_read :  STD_LOGIC;
                signal analyzer_input_left_avalon_slave_readdata :  STD_LOGIC_VECTOR (127 DOWNTO 0);
                signal analyzer_input_left_avalon_slave_readdata_from_sa :  STD_LOGIC_VECTOR (127 DOWNTO 0);
                signal analyzer_input_left_avalon_slave_reset_n :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_read :  STD_LOGIC;
                signal analyzer_input_right_avalon_slave_readdata :  STD_LOGIC_VECTOR (127 DOWNTO 0);
                signal analyzer_input_right_avalon_slave_readdata_from_sa :  STD_LOGIC_VECTOR (127 DOWNTO 0);
                signal analyzer_input_right_avalon_slave_reset_n :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal audio_and_video_config_0_avalon_on_board_config_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal audio_and_video_config_0_avalon_on_board_config_slave_chipselect :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_read :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal audio_and_video_config_0_avalon_on_board_config_slave_reset :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_write :  STD_LOGIC;
                signal audio_and_video_config_0_avalon_on_board_config_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal character_buffer_avalon_char_buffer_slave_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal character_buffer_avalon_char_buffer_slave_chipselect :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_read :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal character_buffer_avalon_char_buffer_slave_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal character_buffer_avalon_char_buffer_slave_waitrequest :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_waitrequest_from_sa :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_write :  STD_LOGIC;
                signal character_buffer_avalon_char_buffer_slave_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal character_buffer_avalon_char_control_slave_address :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal character_buffer_avalon_char_control_slave_chipselect :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_read :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal character_buffer_avalon_char_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal character_buffer_avalon_char_control_slave_reset :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_write :  STD_LOGIC;
                signal character_buffer_avalon_char_control_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal character_buffer_avalon_char_source_data :  STD_LOGIC_VECTOR (39 DOWNTO 0);
                signal character_buffer_avalon_char_source_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal character_buffer_avalon_char_source_endofpacket :  STD_LOGIC;
                signal character_buffer_avalon_char_source_ready :  STD_LOGIC;
                signal character_buffer_avalon_char_source_startofpacket :  STD_LOGIC;
                signal character_buffer_avalon_char_source_valid :  STD_LOGIC;
                signal clk_0_reset_n :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_clk_en :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_done :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_estatus :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_n :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_readra :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_readrb :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_start :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_status :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_writerc :  STD_LOGIC;
                signal cpu_custom_instruction_master_reset_n :  STD_LOGIC;
                signal cpu_custom_instruction_master_start_cpu_fpoint_s1 :  STD_LOGIC;
                signal cpu_data_master_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_byteenable_sdram_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_byteenable_sram_avalon_sram_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_data_master_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal cpu_data_master_dbs_write_8 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal cpu_data_master_debugaccess :  STD_LOGIC;
                signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal cpu_data_master_granted_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_granted_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal cpu_data_master_granted_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_granted_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal cpu_data_master_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_data_master_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpu_data_master_granted_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_compressor_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_delay_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_delay_decay_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_delay_length_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_master_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_output_power_left_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_output_power_right_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_granted_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal cpu_data_master_granted_sdram_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_data_master_no_byte_enables_and_last_term :  STD_LOGIC;
                signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal cpu_data_master_qualified_request_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_compressor_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_delay_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_delay_decay_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_delay_length_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_master_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_output_power_left_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_output_power_right_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal cpu_data_master_qualified_request_sdram_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_data_master_read :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_compressor_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_delay_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_delay_decay_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_delay_length_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_master_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_output_power_left_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_output_power_right_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data :  STD_LOGIC;
                signal cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control :  STD_LOGIC;
                signal cpu_data_master_requests_analyzer_input_left_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_requests_analyzer_input_right_avalon_slave :  STD_LOGIC;
                signal cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal cpu_data_master_requests_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_requests_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal cpu_data_master_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_data_master_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpu_data_master_requests_pio_bitcrusher_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_bitcrusher_crush_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_bitcrusher_downsample_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_bitcrusher_drywet_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_bitcrusher_flavor_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_bitcrusher_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_compressor_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_compressor_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_compressor_treshold_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_delay_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_delay_decay_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_delay_length_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_master_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_octaver_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_octaver_dry_wet_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_output_power_left_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_output_power_right_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_overdrive_asymmetric_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_overdrive_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_overdrive_gain_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_overdrive_tone_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_overdrive_volume_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_tremolo_stereo_depth_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_tremolo_stereo_mode_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal cpu_data_master_requests_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal cpu_data_master_requests_sdram_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_data_master_waitrequest :  STD_LOGIC;
                signal cpu_data_master_write :  STD_LOGIC;
                signal cpu_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_fpoint_s1_clk_en :  STD_LOGIC;
                signal cpu_fpoint_s1_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_fpoint_s1_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_fpoint_s1_done :  STD_LOGIC;
                signal cpu_fpoint_s1_done_from_sa :  STD_LOGIC;
                signal cpu_fpoint_s1_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_fpoint_s1_reset :  STD_LOGIC;
                signal cpu_fpoint_s1_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_fpoint_s1_result_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_fpoint_s1_select :  STD_LOGIC;
                signal cpu_fpoint_s1_start :  STD_LOGIC;
                signal cpu_instruction_master_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_instruction_master_granted_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_instruction_master_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_instruction_master_read :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal cpu_instruction_master_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal cpu_instruction_master_requests_sram_avalon_sram_slave :  STD_LOGIC;
                signal cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal cpu_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_chipselect :  STD_LOGIC;
                signal cpu_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal cpu_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal cpu_jtag_debug_module_write :  STD_LOGIC;
                signal cpu_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer :  STD_LOGIC;
                signal d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer :  STD_LOGIC;
                signal d1_analyzer_input_left_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_analyzer_input_right_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer :  STD_LOGIC;
                signal d1_character_buffer_avalon_char_buffer_slave_end_xfer :  STD_LOGIC;
                signal d1_character_buffer_avalon_char_control_slave_end_xfer :  STD_LOGIC;
                signal d1_cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_pio_bitcrusher_bypass_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_bitcrusher_crush_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_bitcrusher_downsample_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_bitcrusher_drywet_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_bitcrusher_flavor_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_bitcrusher_tone_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_compressor_bypass_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_compressor_gain_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_compressor_treshold_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_delay_bypass_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_delay_decay_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_delay_length_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_master_volume_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_octaver_bypass_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_octaver_dry_wet_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_output_power_left_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_output_power_right_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_overdrive_asymmetric_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_overdrive_bypass_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_overdrive_gain_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_overdrive_tone_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_overdrive_volume_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_tremolo_stereo_bypass_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_tremolo_stereo_depth_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_tremolo_stereo_mode_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_tremolo_stereo_sweep_a_s1_end_xfer :  STD_LOGIC;
                signal d1_pio_tremolo_stereo_sweep_b_s1_end_xfer :  STD_LOGIC;
                signal d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer :  STD_LOGIC;
                signal d1_ps2_avalon_ps2_slave_end_xfer :  STD_LOGIC;
                signal d1_sdram_s1_end_xfer :  STD_LOGIC;
                signal d1_sram_avalon_sram_slave_end_xfer :  STD_LOGIC;
                signal internal_FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal internal_FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal internal_FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal internal_FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal internal_FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal internal_I2C_SCLK_from_the_audio_and_video_config_0 :  STD_LOGIC;
                signal internal_SRAM_ADDR_from_the_sram :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal internal_SRAM_CE_N_from_the_sram :  STD_LOGIC;
                signal internal_SRAM_LB_N_from_the_sram :  STD_LOGIC;
                signal internal_SRAM_OE_N_from_the_sram :  STD_LOGIC;
                signal internal_SRAM_UB_N_from_the_sram :  STD_LOGIC;
                signal internal_SRAM_WE_N_from_the_sram :  STD_LOGIC;
                signal internal_VGA_BLANK_from_the_vga :  STD_LOGIC;
                signal internal_VGA_B_from_the_vga :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_VGA_G_from_the_vga :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_VGA_HS_from_the_vga :  STD_LOGIC;
                signal internal_VGA_R_from_the_vga :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_VGA_SYNC_from_the_vga :  STD_LOGIC;
                signal internal_VGA_VS_from_the_vga :  STD_LOGIC;
                signal internal_out_port_from_the_pio_bitcrusher_bypass :  STD_LOGIC;
                signal internal_out_port_from_the_pio_bitcrusher_crush :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_out_port_from_the_pio_bitcrusher_downsample :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_pio_bitcrusher_drywet :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_bitcrusher_flavor :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_out_port_from_the_pio_bitcrusher_tone :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_compressor_bypass :  STD_LOGIC;
                signal internal_out_port_from_the_pio_compressor_gain :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_pio_compressor_treshold :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_delay_bypass :  STD_LOGIC;
                signal internal_out_port_from_the_pio_delay_decay :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_pio_delay_length :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_master_volume :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_octaver_bypass :  STD_LOGIC;
                signal internal_out_port_from_the_pio_octaver_dry_wet :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_overdrive_asymmetric :  STD_LOGIC;
                signal internal_out_port_from_the_pio_overdrive_bypass :  STD_LOGIC;
                signal internal_out_port_from_the_pio_overdrive_gain :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_overdrive_tone :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_overdrive_volume :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_tremolo_stereo_bypass :  STD_LOGIC;
                signal internal_out_port_from_the_pio_tremolo_stereo_depth :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_out_port_from_the_pio_tremolo_stereo_mode :  STD_LOGIC;
                signal internal_out_port_from_the_pio_tremolo_stereo_sweep_a :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_out_port_from_the_pio_tremolo_stereo_sweep_b :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_sample_left_out_from_the_membuffer_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_sample_right_out_from_the_membuffer_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_zs_addr_from_the_sdram :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal internal_zs_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_cas_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_cke_from_the_sdram :  STD_LOGIC;
                signal internal_zs_cs_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_dqm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_ras_n_from_the_sdram :  STD_LOGIC;
                signal internal_zs_we_n_from_the_sdram :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal membuffer_0_avalon_master_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal membuffer_0_avalon_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal membuffer_0_avalon_master_read :  STD_LOGIC;
                signal membuffer_0_avalon_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal membuffer_0_avalon_master_reset_n :  STD_LOGIC;
                signal membuffer_0_avalon_master_waitrequest :  STD_LOGIC;
                signal membuffer_0_avalon_master_write :  STD_LOGIC;
                signal membuffer_0_avalon_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal membuffer_0_byteenable_sdram_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal membuffer_0_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal membuffer_0_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal membuffer_0_granted_sdram_s1 :  STD_LOGIC;
                signal membuffer_0_qualified_request_sdram_s1 :  STD_LOGIC;
                signal membuffer_0_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal membuffer_0_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal membuffer_0_requests_sdram_s1 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_bitcrusher_bypass_s1_chipselect :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_readdata :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_reset_n :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_write_n :  STD_LOGIC;
                signal pio_bitcrusher_bypass_s1_writedata :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_bitcrusher_crush_s1_chipselect :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_readdata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_bitcrusher_crush_s1_readdata_from_sa :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_bitcrusher_crush_s1_reset_n :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_write_n :  STD_LOGIC;
                signal pio_bitcrusher_crush_s1_writedata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_bitcrusher_downsample_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_bitcrusher_downsample_s1_chipselect :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_bitcrusher_downsample_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_bitcrusher_downsample_s1_reset_n :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_write_n :  STD_LOGIC;
                signal pio_bitcrusher_downsample_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_bitcrusher_drywet_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_bitcrusher_drywet_s1_chipselect :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_bitcrusher_drywet_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_bitcrusher_drywet_s1_reset_n :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_write_n :  STD_LOGIC;
                signal pio_bitcrusher_drywet_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_bitcrusher_flavor_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_bitcrusher_flavor_s1_chipselect :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_readdata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_bitcrusher_flavor_s1_readdata_from_sa :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_bitcrusher_flavor_s1_reset_n :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_write_n :  STD_LOGIC;
                signal pio_bitcrusher_flavor_s1_writedata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_bitcrusher_tone_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_bitcrusher_tone_s1_chipselect :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_bitcrusher_tone_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_bitcrusher_tone_s1_reset_n :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_write_n :  STD_LOGIC;
                signal pio_bitcrusher_tone_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_compressor_bypass_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_compressor_bypass_s1_chipselect :  STD_LOGIC;
                signal pio_compressor_bypass_s1_readdata :  STD_LOGIC;
                signal pio_compressor_bypass_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_compressor_bypass_s1_reset_n :  STD_LOGIC;
                signal pio_compressor_bypass_s1_write_n :  STD_LOGIC;
                signal pio_compressor_bypass_s1_writedata :  STD_LOGIC;
                signal pio_compressor_gain_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_compressor_gain_s1_chipselect :  STD_LOGIC;
                signal pio_compressor_gain_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_compressor_gain_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_compressor_gain_s1_reset_n :  STD_LOGIC;
                signal pio_compressor_gain_s1_write_n :  STD_LOGIC;
                signal pio_compressor_gain_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_compressor_treshold_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_compressor_treshold_s1_chipselect :  STD_LOGIC;
                signal pio_compressor_treshold_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_compressor_treshold_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_compressor_treshold_s1_reset_n :  STD_LOGIC;
                signal pio_compressor_treshold_s1_write_n :  STD_LOGIC;
                signal pio_compressor_treshold_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_delay_bypass_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_delay_bypass_s1_chipselect :  STD_LOGIC;
                signal pio_delay_bypass_s1_readdata :  STD_LOGIC;
                signal pio_delay_bypass_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_delay_bypass_s1_reset_n :  STD_LOGIC;
                signal pio_delay_bypass_s1_write_n :  STD_LOGIC;
                signal pio_delay_bypass_s1_writedata :  STD_LOGIC;
                signal pio_delay_decay_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_delay_decay_s1_chipselect :  STD_LOGIC;
                signal pio_delay_decay_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_delay_decay_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_delay_decay_s1_reset_n :  STD_LOGIC;
                signal pio_delay_decay_s1_write_n :  STD_LOGIC;
                signal pio_delay_decay_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pio_delay_length_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_delay_length_s1_chipselect :  STD_LOGIC;
                signal pio_delay_length_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_delay_length_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_delay_length_s1_reset_n :  STD_LOGIC;
                signal pio_delay_length_s1_write_n :  STD_LOGIC;
                signal pio_delay_length_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_master_volume_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_master_volume_s1_chipselect :  STD_LOGIC;
                signal pio_master_volume_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_master_volume_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_master_volume_s1_reset_n :  STD_LOGIC;
                signal pio_master_volume_s1_write_n :  STD_LOGIC;
                signal pio_master_volume_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_octaver_bypass_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_octaver_bypass_s1_chipselect :  STD_LOGIC;
                signal pio_octaver_bypass_s1_readdata :  STD_LOGIC;
                signal pio_octaver_bypass_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_octaver_bypass_s1_reset_n :  STD_LOGIC;
                signal pio_octaver_bypass_s1_write_n :  STD_LOGIC;
                signal pio_octaver_bypass_s1_writedata :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_octaver_dry_wet_s1_chipselect :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_octaver_dry_wet_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_octaver_dry_wet_s1_reset_n :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_write_n :  STD_LOGIC;
                signal pio_octaver_dry_wet_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_output_power_left_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_output_power_left_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_output_power_left_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_output_power_left_s1_reset_n :  STD_LOGIC;
                signal pio_output_power_right_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_output_power_right_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_output_power_right_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_output_power_right_s1_reset_n :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_overdrive_asymmetric_s1_chipselect :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_readdata :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_reset_n :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_write_n :  STD_LOGIC;
                signal pio_overdrive_asymmetric_s1_writedata :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_overdrive_bypass_s1_chipselect :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_readdata :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_reset_n :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_write_n :  STD_LOGIC;
                signal pio_overdrive_bypass_s1_writedata :  STD_LOGIC;
                signal pio_overdrive_gain_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_overdrive_gain_s1_chipselect :  STD_LOGIC;
                signal pio_overdrive_gain_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_gain_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_gain_s1_reset_n :  STD_LOGIC;
                signal pio_overdrive_gain_s1_write_n :  STD_LOGIC;
                signal pio_overdrive_gain_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_tone_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_overdrive_tone_s1_chipselect :  STD_LOGIC;
                signal pio_overdrive_tone_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_tone_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_tone_s1_reset_n :  STD_LOGIC;
                signal pio_overdrive_tone_s1_write_n :  STD_LOGIC;
                signal pio_overdrive_tone_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_volume_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_overdrive_volume_s1_chipselect :  STD_LOGIC;
                signal pio_overdrive_volume_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_volume_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_overdrive_volume_s1_reset_n :  STD_LOGIC;
                signal pio_overdrive_volume_s1_write_n :  STD_LOGIC;
                signal pio_overdrive_volume_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_tremolo_stereo_bypass_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_tremolo_stereo_bypass_s1_chipselect :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_readdata :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_reset_n :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_write_n :  STD_LOGIC;
                signal pio_tremolo_stereo_bypass_s1_writedata :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_tremolo_stereo_depth_s1_chipselect :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_tremolo_stereo_depth_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_tremolo_stereo_depth_s1_reset_n :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_write_n :  STD_LOGIC;
                signal pio_tremolo_stereo_depth_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pio_tremolo_stereo_mode_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_tremolo_stereo_mode_s1_chipselect :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_readdata :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_readdata_from_sa :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_reset_n :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_write_n :  STD_LOGIC;
                signal pio_tremolo_stereo_mode_s1_writedata :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_a_s1_chipselect :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_readdata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_a_s1_readdata_from_sa :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_a_s1_reset_n :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_write_n :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_a_s1_writedata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_b_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_b_s1_chipselect :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_readdata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_b_s1_readdata_from_sa :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pio_tremolo_stereo_sweep_b_s1_reset_n :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_write_n :  STD_LOGIC;
                signal pio_tremolo_stereo_sweep_b_s1_writedata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_master_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_master_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_master_arbiterlock :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_latency_counter :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_read :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_master_readdatavalid :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_master_waitrequest :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_slave_read :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_slave_reset :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_write :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_source_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_source_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pixel_buffer_avalon_pixel_buffer_source_endofpacket :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_source_ready :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_source_startofpacket :  STD_LOGIC;
                signal pixel_buffer_avalon_pixel_buffer_source_valid :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_address :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ps2_avalon_ps2_slave_chipselect :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_irq :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_irq_from_sa :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_read :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ps2_avalon_ps2_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ps2_avalon_ps2_slave_reset :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_waitrequest :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_waitrequest_from_sa :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_write :  STD_LOGIC;
                signal ps2_avalon_ps2_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave :  STD_LOGIC;
                signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave :  STD_LOGIC;
                signal registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave :  STD_LOGIC;
                signal registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave :  STD_LOGIC;
                signal registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave :  STD_LOGIC;
                signal registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave :  STD_LOGIC;
                signal reset_n_sources :  STD_LOGIC;
                signal sdram_s1_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal sdram_s1_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_s1_chipselect :  STD_LOGIC;
                signal sdram_s1_read_n :  STD_LOGIC;
                signal sdram_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sdram_s1_readdatavalid :  STD_LOGIC;
                signal sdram_s1_reset_n :  STD_LOGIC;
                signal sdram_s1_waitrequest :  STD_LOGIC;
                signal sdram_s1_waitrequest_from_sa :  STD_LOGIC;
                signal sdram_s1_write_n :  STD_LOGIC;
                signal sdram_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sram_avalon_sram_slave_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal sram_avalon_sram_slave_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sram_avalon_sram_slave_read :  STD_LOGIC;
                signal sram_avalon_sram_slave_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sram_avalon_sram_slave_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sram_avalon_sram_slave_reset :  STD_LOGIC;
                signal sram_avalon_sram_slave_write :  STD_LOGIC;
                signal sram_avalon_sram_slave_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal vga_avalon_vga_sink_data :  STD_LOGIC_VECTOR (29 DOWNTO 0);
                signal vga_avalon_vga_sink_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal vga_avalon_vga_sink_endofpacket :  STD_LOGIC;
                signal vga_avalon_vga_sink_ready :  STD_LOGIC;
                signal vga_avalon_vga_sink_ready_from_sa :  STD_LOGIC;
                signal vga_avalon_vga_sink_reset :  STD_LOGIC;
                signal vga_avalon_vga_sink_startofpacket :  STD_LOGIC;
                signal vga_avalon_vga_sink_valid :  STD_LOGIC;

begin

  --the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data, which is an e_instance
  the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data : Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_arbitrator
    port map(
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata,
      cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer => d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      reset_n => clk_0_reset_n
    );


  --the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control, which is an e_instance
  the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control : Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_arbitrator
    port map(
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata,
      cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer => d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      reset_n => clk_0_reset_n
    );


  --the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0, which is an e_ptf_instance
  the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0
    port map(
      FL_ADDR => internal_FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_CE_N => internal_FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_DQ => FL_DQ_to_and_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_OE_N => internal_FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_RST_N => internal_FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_WE_N => internal_FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      o_avalon_erase_readdata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata,
      o_avalon_erase_waitrequest => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest,
      o_avalon_readdata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata,
      o_avalon_waitrequest => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest,
      i_avalon_address => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address,
      i_avalon_byteenable => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable,
      i_avalon_chip_select => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect,
      i_avalon_erase_byteenable => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable,
      i_avalon_erase_chip_select => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect,
      i_avalon_erase_read => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read,
      i_avalon_erase_write => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write,
      i_avalon_erase_writedata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata,
      i_avalon_read => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read,
      i_avalon_write => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write,
      i_avalon_writedata => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata,
      i_clock => clk_0,
      i_reset_n => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_reset_n
    );


  --the_alpha_blending_avalon_background_sink, which is an e_instance
  the_alpha_blending_avalon_background_sink : alpha_blending_avalon_background_sink_arbitrator
    port map(
      alpha_blending_avalon_background_sink_data => alpha_blending_avalon_background_sink_data,
      alpha_blending_avalon_background_sink_empty => alpha_blending_avalon_background_sink_empty,
      alpha_blending_avalon_background_sink_endofpacket => alpha_blending_avalon_background_sink_endofpacket,
      alpha_blending_avalon_background_sink_ready_from_sa => alpha_blending_avalon_background_sink_ready_from_sa,
      alpha_blending_avalon_background_sink_startofpacket => alpha_blending_avalon_background_sink_startofpacket,
      alpha_blending_avalon_background_sink_valid => alpha_blending_avalon_background_sink_valid,
      alpha_blending_avalon_background_sink_ready => alpha_blending_avalon_background_sink_ready,
      clk => clk_0,
      pixel_buffer_avalon_pixel_buffer_source_data => pixel_buffer_avalon_pixel_buffer_source_data,
      pixel_buffer_avalon_pixel_buffer_source_empty => pixel_buffer_avalon_pixel_buffer_source_empty,
      pixel_buffer_avalon_pixel_buffer_source_endofpacket => pixel_buffer_avalon_pixel_buffer_source_endofpacket,
      pixel_buffer_avalon_pixel_buffer_source_startofpacket => pixel_buffer_avalon_pixel_buffer_source_startofpacket,
      pixel_buffer_avalon_pixel_buffer_source_valid => pixel_buffer_avalon_pixel_buffer_source_valid,
      reset_n => clk_0_reset_n
    );


  --the_alpha_blending_avalon_foreground_sink, which is an e_instance
  the_alpha_blending_avalon_foreground_sink : alpha_blending_avalon_foreground_sink_arbitrator
    port map(
      alpha_blending_avalon_foreground_sink_data => alpha_blending_avalon_foreground_sink_data,
      alpha_blending_avalon_foreground_sink_empty => alpha_blending_avalon_foreground_sink_empty,
      alpha_blending_avalon_foreground_sink_endofpacket => alpha_blending_avalon_foreground_sink_endofpacket,
      alpha_blending_avalon_foreground_sink_ready_from_sa => alpha_blending_avalon_foreground_sink_ready_from_sa,
      alpha_blending_avalon_foreground_sink_reset => alpha_blending_avalon_foreground_sink_reset,
      alpha_blending_avalon_foreground_sink_startofpacket => alpha_blending_avalon_foreground_sink_startofpacket,
      alpha_blending_avalon_foreground_sink_valid => alpha_blending_avalon_foreground_sink_valid,
      alpha_blending_avalon_foreground_sink_ready => alpha_blending_avalon_foreground_sink_ready,
      character_buffer_avalon_char_source_data => character_buffer_avalon_char_source_data,
      character_buffer_avalon_char_source_empty => character_buffer_avalon_char_source_empty,
      character_buffer_avalon_char_source_endofpacket => character_buffer_avalon_char_source_endofpacket,
      character_buffer_avalon_char_source_startofpacket => character_buffer_avalon_char_source_startofpacket,
      character_buffer_avalon_char_source_valid => character_buffer_avalon_char_source_valid,
      clk => clk_0,
      reset_n => clk_0_reset_n
    );


  --the_alpha_blending_avalon_blended_source, which is an e_instance
  the_alpha_blending_avalon_blended_source : alpha_blending_avalon_blended_source_arbitrator
    port map(
      alpha_blending_avalon_blended_source_ready => alpha_blending_avalon_blended_source_ready,
      alpha_blending_avalon_blended_source_data => alpha_blending_avalon_blended_source_data,
      alpha_blending_avalon_blended_source_empty => alpha_blending_avalon_blended_source_empty,
      alpha_blending_avalon_blended_source_endofpacket => alpha_blending_avalon_blended_source_endofpacket,
      alpha_blending_avalon_blended_source_startofpacket => alpha_blending_avalon_blended_source_startofpacket,
      alpha_blending_avalon_blended_source_valid => alpha_blending_avalon_blended_source_valid,
      clk => clk_0,
      reset_n => clk_0_reset_n,
      vga_avalon_vga_sink_ready_from_sa => vga_avalon_vga_sink_ready_from_sa
    );


  --the_alpha_blending, which is an e_ptf_instance
  the_alpha_blending : alpha_blending
    port map(
      background_ready => alpha_blending_avalon_background_sink_ready,
      foreground_ready => alpha_blending_avalon_foreground_sink_ready,
      output_data => alpha_blending_avalon_blended_source_data,
      output_empty => alpha_blending_avalon_blended_source_empty,
      output_endofpacket => alpha_blending_avalon_blended_source_endofpacket,
      output_startofpacket => alpha_blending_avalon_blended_source_startofpacket,
      output_valid => alpha_blending_avalon_blended_source_valid,
      background_data => alpha_blending_avalon_background_sink_data,
      background_empty => alpha_blending_avalon_background_sink_empty,
      background_endofpacket => alpha_blending_avalon_background_sink_endofpacket,
      background_startofpacket => alpha_blending_avalon_background_sink_startofpacket,
      background_valid => alpha_blending_avalon_background_sink_valid,
      clk => clk_0,
      foreground_data => alpha_blending_avalon_foreground_sink_data,
      foreground_empty => alpha_blending_avalon_foreground_sink_empty,
      foreground_endofpacket => alpha_blending_avalon_foreground_sink_endofpacket,
      foreground_startofpacket => alpha_blending_avalon_foreground_sink_startofpacket,
      foreground_valid => alpha_blending_avalon_foreground_sink_valid,
      output_ready => alpha_blending_avalon_blended_source_ready,
      reset => alpha_blending_avalon_foreground_sink_reset
    );


  --the_analyzer_input_left_avalon_slave, which is an e_instance
  the_analyzer_input_left_avalon_slave : analyzer_input_left_avalon_slave_arbitrator
    port map(
      analyzer_input_left_avalon_slave_read => analyzer_input_left_avalon_slave_read,
      analyzer_input_left_avalon_slave_readdata_from_sa => analyzer_input_left_avalon_slave_readdata_from_sa,
      analyzer_input_left_avalon_slave_reset_n => analyzer_input_left_avalon_slave_reset_n,
      cpu_data_master_granted_analyzer_input_left_avalon_slave => cpu_data_master_granted_analyzer_input_left_avalon_slave,
      cpu_data_master_qualified_request_analyzer_input_left_avalon_slave => cpu_data_master_qualified_request_analyzer_input_left_avalon_slave,
      cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave => cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave,
      cpu_data_master_requests_analyzer_input_left_avalon_slave => cpu_data_master_requests_analyzer_input_left_avalon_slave,
      d1_analyzer_input_left_avalon_slave_end_xfer => d1_analyzer_input_left_avalon_slave_end_xfer,
      analyzer_input_left_avalon_slave_readdata => analyzer_input_left_avalon_slave_readdata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_write => cpu_data_master_write,
      reset_n => clk_0_reset_n
    );


  --the_analyzer_input_left, which is an e_ptf_instance
  the_analyzer_input_left : analyzer_input_left
    port map(
      readdata => analyzer_input_left_avalon_slave_readdata,
      clk => clk_0,
      read => analyzer_input_left_avalon_slave_read,
      reset => analyzer_input_left_avalon_slave_reset_n,
      x_in => x_in_to_the_analyzer_input_left,
      y_in => y_in_to_the_analyzer_input_left
    );


  --the_analyzer_input_right_avalon_slave, which is an e_instance
  the_analyzer_input_right_avalon_slave : analyzer_input_right_avalon_slave_arbitrator
    port map(
      analyzer_input_right_avalon_slave_read => analyzer_input_right_avalon_slave_read,
      analyzer_input_right_avalon_slave_readdata_from_sa => analyzer_input_right_avalon_slave_readdata_from_sa,
      analyzer_input_right_avalon_slave_reset_n => analyzer_input_right_avalon_slave_reset_n,
      cpu_data_master_granted_analyzer_input_right_avalon_slave => cpu_data_master_granted_analyzer_input_right_avalon_slave,
      cpu_data_master_qualified_request_analyzer_input_right_avalon_slave => cpu_data_master_qualified_request_analyzer_input_right_avalon_slave,
      cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave => cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave,
      cpu_data_master_requests_analyzer_input_right_avalon_slave => cpu_data_master_requests_analyzer_input_right_avalon_slave,
      d1_analyzer_input_right_avalon_slave_end_xfer => d1_analyzer_input_right_avalon_slave_end_xfer,
      analyzer_input_right_avalon_slave_readdata => analyzer_input_right_avalon_slave_readdata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_write => cpu_data_master_write,
      reset_n => clk_0_reset_n
    );


  --the_analyzer_input_right, which is an e_ptf_instance
  the_analyzer_input_right : analyzer_input_right
    port map(
      readdata => analyzer_input_right_avalon_slave_readdata,
      clk => clk_0,
      read => analyzer_input_right_avalon_slave_read,
      reset => analyzer_input_right_avalon_slave_reset_n,
      x_in => x_in_to_the_analyzer_input_right,
      y_in => y_in_to_the_analyzer_input_right
    );


  --the_audio_and_video_config_0_avalon_on_board_config_slave, which is an e_instance
  the_audio_and_video_config_0_avalon_on_board_config_slave : audio_and_video_config_0_avalon_on_board_config_slave_arbitrator
    port map(
      audio_and_video_config_0_avalon_on_board_config_slave_address => audio_and_video_config_0_avalon_on_board_config_slave_address,
      audio_and_video_config_0_avalon_on_board_config_slave_byteenable => audio_and_video_config_0_avalon_on_board_config_slave_byteenable,
      audio_and_video_config_0_avalon_on_board_config_slave_chipselect => audio_and_video_config_0_avalon_on_board_config_slave_chipselect,
      audio_and_video_config_0_avalon_on_board_config_slave_read => audio_and_video_config_0_avalon_on_board_config_slave_read,
      audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa => audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa,
      audio_and_video_config_0_avalon_on_board_config_slave_reset => audio_and_video_config_0_avalon_on_board_config_slave_reset,
      audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa => audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa,
      audio_and_video_config_0_avalon_on_board_config_slave_write => audio_and_video_config_0_avalon_on_board_config_slave_write,
      audio_and_video_config_0_avalon_on_board_config_slave_writedata => audio_and_video_config_0_avalon_on_board_config_slave_writedata,
      cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave,
      cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave,
      cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave,
      cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave,
      d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer => d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer,
      registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave => registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave,
      audio_and_video_config_0_avalon_on_board_config_slave_readdata => audio_and_video_config_0_avalon_on_board_config_slave_readdata,
      audio_and_video_config_0_avalon_on_board_config_slave_waitrequest => audio_and_video_config_0_avalon_on_board_config_slave_waitrequest,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      reset_n => clk_0_reset_n
    );


  --the_audio_and_video_config_0, which is an e_ptf_instance
  the_audio_and_video_config_0 : audio_and_video_config_0
    port map(
      I2C_SCLK => internal_I2C_SCLK_from_the_audio_and_video_config_0,
      I2C_SDAT => I2C_SDAT_to_and_from_the_audio_and_video_config_0,
      ob_readdata => audio_and_video_config_0_avalon_on_board_config_slave_readdata,
      ob_waitrequest => audio_and_video_config_0_avalon_on_board_config_slave_waitrequest,
      clk => clk_0,
      ob_address => audio_and_video_config_0_avalon_on_board_config_slave_address,
      ob_byteenable => audio_and_video_config_0_avalon_on_board_config_slave_byteenable,
      ob_chipselect => audio_and_video_config_0_avalon_on_board_config_slave_chipselect,
      ob_read => audio_and_video_config_0_avalon_on_board_config_slave_read,
      ob_write => audio_and_video_config_0_avalon_on_board_config_slave_write,
      ob_writedata => audio_and_video_config_0_avalon_on_board_config_slave_writedata,
      reset => audio_and_video_config_0_avalon_on_board_config_slave_reset
    );


  --the_character_buffer_avalon_char_buffer_slave, which is an e_instance
  the_character_buffer_avalon_char_buffer_slave : character_buffer_avalon_char_buffer_slave_arbitrator
    port map(
      character_buffer_avalon_char_buffer_slave_address => character_buffer_avalon_char_buffer_slave_address,
      character_buffer_avalon_char_buffer_slave_chipselect => character_buffer_avalon_char_buffer_slave_chipselect,
      character_buffer_avalon_char_buffer_slave_read => character_buffer_avalon_char_buffer_slave_read,
      character_buffer_avalon_char_buffer_slave_readdata_from_sa => character_buffer_avalon_char_buffer_slave_readdata_from_sa,
      character_buffer_avalon_char_buffer_slave_waitrequest_from_sa => character_buffer_avalon_char_buffer_slave_waitrequest_from_sa,
      character_buffer_avalon_char_buffer_slave_write => character_buffer_avalon_char_buffer_slave_write,
      character_buffer_avalon_char_buffer_slave_writedata => character_buffer_avalon_char_buffer_slave_writedata,
      cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave => cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_granted_character_buffer_avalon_char_buffer_slave => cpu_data_master_granted_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave => cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave => cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_requests_character_buffer_avalon_char_buffer_slave => cpu_data_master_requests_character_buffer_avalon_char_buffer_slave,
      d1_character_buffer_avalon_char_buffer_slave_end_xfer => d1_character_buffer_avalon_char_buffer_slave_end_xfer,
      registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave => registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave,
      character_buffer_avalon_char_buffer_slave_readdata => character_buffer_avalon_char_buffer_slave_readdata,
      character_buffer_avalon_char_buffer_slave_waitrequest => character_buffer_avalon_char_buffer_slave_waitrequest,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_8 => cpu_data_master_dbs_write_8,
      cpu_data_master_no_byte_enables_and_last_term => cpu_data_master_no_byte_enables_and_last_term,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      reset_n => clk_0_reset_n
    );


  --the_character_buffer_avalon_char_control_slave, which is an e_instance
  the_character_buffer_avalon_char_control_slave : character_buffer_avalon_char_control_slave_arbitrator
    port map(
      character_buffer_avalon_char_control_slave_address => character_buffer_avalon_char_control_slave_address,
      character_buffer_avalon_char_control_slave_byteenable => character_buffer_avalon_char_control_slave_byteenable,
      character_buffer_avalon_char_control_slave_chipselect => character_buffer_avalon_char_control_slave_chipselect,
      character_buffer_avalon_char_control_slave_read => character_buffer_avalon_char_control_slave_read,
      character_buffer_avalon_char_control_slave_readdata_from_sa => character_buffer_avalon_char_control_slave_readdata_from_sa,
      character_buffer_avalon_char_control_slave_reset => character_buffer_avalon_char_control_slave_reset,
      character_buffer_avalon_char_control_slave_write => character_buffer_avalon_char_control_slave_write,
      character_buffer_avalon_char_control_slave_writedata => character_buffer_avalon_char_control_slave_writedata,
      cpu_data_master_granted_character_buffer_avalon_char_control_slave => cpu_data_master_granted_character_buffer_avalon_char_control_slave,
      cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave => cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave,
      cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave => cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave,
      cpu_data_master_requests_character_buffer_avalon_char_control_slave => cpu_data_master_requests_character_buffer_avalon_char_control_slave,
      d1_character_buffer_avalon_char_control_slave_end_xfer => d1_character_buffer_avalon_char_control_slave_end_xfer,
      registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave => registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave,
      character_buffer_avalon_char_control_slave_readdata => character_buffer_avalon_char_control_slave_readdata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      reset_n => clk_0_reset_n
    );


  --the_character_buffer_avalon_char_source, which is an e_instance
  the_character_buffer_avalon_char_source : character_buffer_avalon_char_source_arbitrator
    port map(
      character_buffer_avalon_char_source_ready => character_buffer_avalon_char_source_ready,
      alpha_blending_avalon_foreground_sink_ready_from_sa => alpha_blending_avalon_foreground_sink_ready_from_sa,
      character_buffer_avalon_char_source_data => character_buffer_avalon_char_source_data,
      character_buffer_avalon_char_source_empty => character_buffer_avalon_char_source_empty,
      character_buffer_avalon_char_source_endofpacket => character_buffer_avalon_char_source_endofpacket,
      character_buffer_avalon_char_source_startofpacket => character_buffer_avalon_char_source_startofpacket,
      character_buffer_avalon_char_source_valid => character_buffer_avalon_char_source_valid,
      clk => clk_0,
      reset_n => clk_0_reset_n
    );


  --the_character_buffer, which is an e_ptf_instance
  the_character_buffer : character_buffer
    port map(
      buf_readdata => character_buffer_avalon_char_buffer_slave_readdata,
      buf_waitrequest => character_buffer_avalon_char_buffer_slave_waitrequest,
      ctrl_readdata => character_buffer_avalon_char_control_slave_readdata,
      stream_data => character_buffer_avalon_char_source_data,
      stream_empty => character_buffer_avalon_char_source_empty,
      stream_endofpacket => character_buffer_avalon_char_source_endofpacket,
      stream_startofpacket => character_buffer_avalon_char_source_startofpacket,
      stream_valid => character_buffer_avalon_char_source_valid,
      buf_address => character_buffer_avalon_char_buffer_slave_address,
      buf_chipselect => character_buffer_avalon_char_buffer_slave_chipselect,
      buf_read => character_buffer_avalon_char_buffer_slave_read,
      buf_write => character_buffer_avalon_char_buffer_slave_write,
      buf_writedata => character_buffer_avalon_char_buffer_slave_writedata,
      clk => clk_0,
      ctrl_address => character_buffer_avalon_char_control_slave_address,
      ctrl_byteenable => character_buffer_avalon_char_control_slave_byteenable,
      ctrl_chipselect => character_buffer_avalon_char_control_slave_chipselect,
      ctrl_read => character_buffer_avalon_char_control_slave_read,
      ctrl_write => character_buffer_avalon_char_control_slave_write,
      ctrl_writedata => character_buffer_avalon_char_control_slave_writedata,
      reset => character_buffer_avalon_char_control_slave_reset,
      stream_ready => character_buffer_avalon_char_source_ready
    );


  --the_cpu_jtag_debug_module, which is an e_instance
  the_cpu_jtag_debug_module : cpu_jtag_debug_module_arbitrator
    port map(
      cpu_data_master_granted_cpu_jtag_debug_module => cpu_data_master_granted_cpu_jtag_debug_module,
      cpu_data_master_qualified_request_cpu_jtag_debug_module => cpu_data_master_qualified_request_cpu_jtag_debug_module,
      cpu_data_master_read_data_valid_cpu_jtag_debug_module => cpu_data_master_read_data_valid_cpu_jtag_debug_module,
      cpu_data_master_requests_cpu_jtag_debug_module => cpu_data_master_requests_cpu_jtag_debug_module,
      cpu_instruction_master_granted_cpu_jtag_debug_module => cpu_instruction_master_granted_cpu_jtag_debug_module,
      cpu_instruction_master_qualified_request_cpu_jtag_debug_module => cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
      cpu_instruction_master_read_data_valid_cpu_jtag_debug_module => cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
      cpu_instruction_master_requests_cpu_jtag_debug_module => cpu_instruction_master_requests_cpu_jtag_debug_module,
      cpu_jtag_debug_module_address => cpu_jtag_debug_module_address,
      cpu_jtag_debug_module_begintransfer => cpu_jtag_debug_module_begintransfer,
      cpu_jtag_debug_module_byteenable => cpu_jtag_debug_module_byteenable,
      cpu_jtag_debug_module_chipselect => cpu_jtag_debug_module_chipselect,
      cpu_jtag_debug_module_debugaccess => cpu_jtag_debug_module_debugaccess,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      cpu_jtag_debug_module_resetrequest_from_sa => cpu_jtag_debug_module_resetrequest_from_sa,
      cpu_jtag_debug_module_write => cpu_jtag_debug_module_write,
      cpu_jtag_debug_module_writedata => cpu_jtag_debug_module_writedata,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_jtag_debug_module_readdata => cpu_jtag_debug_module_readdata,
      cpu_jtag_debug_module_resetrequest => cpu_jtag_debug_module_resetrequest,
      reset_n => clk_0_reset_n
    );


  --the_cpu_custom_instruction_master, which is an e_instance
  the_cpu_custom_instruction_master : cpu_custom_instruction_master_arbitrator
    port map(
      cpu_custom_instruction_master_multi_done => cpu_custom_instruction_master_multi_done,
      cpu_custom_instruction_master_multi_result => cpu_custom_instruction_master_multi_result,
      cpu_custom_instruction_master_reset_n => cpu_custom_instruction_master_reset_n,
      cpu_custom_instruction_master_start_cpu_fpoint_s1 => cpu_custom_instruction_master_start_cpu_fpoint_s1,
      cpu_fpoint_s1_select => cpu_fpoint_s1_select,
      clk => clk_0,
      cpu_custom_instruction_master_multi_start => cpu_custom_instruction_master_multi_start,
      cpu_fpoint_s1_done_from_sa => cpu_fpoint_s1_done_from_sa,
      cpu_fpoint_s1_result_from_sa => cpu_fpoint_s1_result_from_sa,
      reset_n => clk_0_reset_n
    );


  --the_cpu_data_master, which is an e_instance
  the_cpu_data_master : cpu_data_master_arbitrator
    port map(
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_16 => cpu_data_master_dbs_write_16,
      cpu_data_master_dbs_write_8 => cpu_data_master_dbs_write_8,
      cpu_data_master_irq => cpu_data_master_irq,
      cpu_data_master_no_byte_enables_and_last_term => cpu_data_master_no_byte_enables_and_last_term,
      cpu_data_master_readdata => cpu_data_master_readdata,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata_from_sa,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest_from_sa,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata_from_sa,
      Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa => Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest_from_sa,
      analyzer_input_left_avalon_slave_readdata_from_sa => analyzer_input_left_avalon_slave_readdata_from_sa,
      analyzer_input_right_avalon_slave_readdata_from_sa => analyzer_input_right_avalon_slave_readdata_from_sa,
      audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa => audio_and_video_config_0_avalon_on_board_config_slave_readdata_from_sa,
      audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa => audio_and_video_config_0_avalon_on_board_config_slave_waitrequest_from_sa,
      character_buffer_avalon_char_buffer_slave_readdata_from_sa => character_buffer_avalon_char_buffer_slave_readdata_from_sa,
      character_buffer_avalon_char_buffer_slave_waitrequest_from_sa => character_buffer_avalon_char_buffer_slave_waitrequest_from_sa,
      character_buffer_avalon_char_control_slave_readdata_from_sa => character_buffer_avalon_char_control_slave_readdata_from_sa,
      clk => clk_0,
      cpu_data_master_address => cpu_data_master_address,
      cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave => cpu_data_master_byteenable_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_byteenable_sdram_s1 => cpu_data_master_byteenable_sdram_s1,
      cpu_data_master_byteenable_sram_avalon_sram_slave => cpu_data_master_byteenable_sram_avalon_sram_slave,
      cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_granted_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      cpu_data_master_granted_analyzer_input_left_avalon_slave => cpu_data_master_granted_analyzer_input_left_avalon_slave,
      cpu_data_master_granted_analyzer_input_right_avalon_slave => cpu_data_master_granted_analyzer_input_right_avalon_slave,
      cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_granted_audio_and_video_config_0_avalon_on_board_config_slave,
      cpu_data_master_granted_character_buffer_avalon_char_buffer_slave => cpu_data_master_granted_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_granted_character_buffer_avalon_char_control_slave => cpu_data_master_granted_character_buffer_avalon_char_control_slave,
      cpu_data_master_granted_cpu_jtag_debug_module => cpu_data_master_granted_cpu_jtag_debug_module,
      cpu_data_master_granted_jtag_uart_avalon_jtag_slave => cpu_data_master_granted_jtag_uart_avalon_jtag_slave,
      cpu_data_master_granted_pio_bitcrusher_bypass_s1 => cpu_data_master_granted_pio_bitcrusher_bypass_s1,
      cpu_data_master_granted_pio_bitcrusher_crush_s1 => cpu_data_master_granted_pio_bitcrusher_crush_s1,
      cpu_data_master_granted_pio_bitcrusher_downsample_s1 => cpu_data_master_granted_pio_bitcrusher_downsample_s1,
      cpu_data_master_granted_pio_bitcrusher_drywet_s1 => cpu_data_master_granted_pio_bitcrusher_drywet_s1,
      cpu_data_master_granted_pio_bitcrusher_flavor_s1 => cpu_data_master_granted_pio_bitcrusher_flavor_s1,
      cpu_data_master_granted_pio_bitcrusher_tone_s1 => cpu_data_master_granted_pio_bitcrusher_tone_s1,
      cpu_data_master_granted_pio_compressor_bypass_s1 => cpu_data_master_granted_pio_compressor_bypass_s1,
      cpu_data_master_granted_pio_compressor_gain_s1 => cpu_data_master_granted_pio_compressor_gain_s1,
      cpu_data_master_granted_pio_compressor_treshold_s1 => cpu_data_master_granted_pio_compressor_treshold_s1,
      cpu_data_master_granted_pio_delay_bypass_s1 => cpu_data_master_granted_pio_delay_bypass_s1,
      cpu_data_master_granted_pio_delay_decay_s1 => cpu_data_master_granted_pio_delay_decay_s1,
      cpu_data_master_granted_pio_delay_length_s1 => cpu_data_master_granted_pio_delay_length_s1,
      cpu_data_master_granted_pio_master_volume_s1 => cpu_data_master_granted_pio_master_volume_s1,
      cpu_data_master_granted_pio_octaver_bypass_s1 => cpu_data_master_granted_pio_octaver_bypass_s1,
      cpu_data_master_granted_pio_octaver_dry_wet_s1 => cpu_data_master_granted_pio_octaver_dry_wet_s1,
      cpu_data_master_granted_pio_output_power_left_s1 => cpu_data_master_granted_pio_output_power_left_s1,
      cpu_data_master_granted_pio_output_power_right_s1 => cpu_data_master_granted_pio_output_power_right_s1,
      cpu_data_master_granted_pio_overdrive_asymmetric_s1 => cpu_data_master_granted_pio_overdrive_asymmetric_s1,
      cpu_data_master_granted_pio_overdrive_bypass_s1 => cpu_data_master_granted_pio_overdrive_bypass_s1,
      cpu_data_master_granted_pio_overdrive_gain_s1 => cpu_data_master_granted_pio_overdrive_gain_s1,
      cpu_data_master_granted_pio_overdrive_tone_s1 => cpu_data_master_granted_pio_overdrive_tone_s1,
      cpu_data_master_granted_pio_overdrive_volume_s1 => cpu_data_master_granted_pio_overdrive_volume_s1,
      cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 => cpu_data_master_granted_pio_tremolo_stereo_bypass_s1,
      cpu_data_master_granted_pio_tremolo_stereo_depth_s1 => cpu_data_master_granted_pio_tremolo_stereo_depth_s1,
      cpu_data_master_granted_pio_tremolo_stereo_mode_s1 => cpu_data_master_granted_pio_tremolo_stereo_mode_s1,
      cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1,
      cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1,
      cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave,
      cpu_data_master_granted_ps2_avalon_ps2_slave => cpu_data_master_granted_ps2_avalon_ps2_slave,
      cpu_data_master_granted_sdram_s1 => cpu_data_master_granted_sdram_s1,
      cpu_data_master_granted_sram_avalon_sram_slave => cpu_data_master_granted_sram_avalon_sram_slave,
      cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_qualified_request_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      cpu_data_master_qualified_request_analyzer_input_left_avalon_slave => cpu_data_master_qualified_request_analyzer_input_left_avalon_slave,
      cpu_data_master_qualified_request_analyzer_input_right_avalon_slave => cpu_data_master_qualified_request_analyzer_input_right_avalon_slave,
      cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_qualified_request_audio_and_video_config_0_avalon_on_board_config_slave,
      cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave => cpu_data_master_qualified_request_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave => cpu_data_master_qualified_request_character_buffer_avalon_char_control_slave,
      cpu_data_master_qualified_request_cpu_jtag_debug_module => cpu_data_master_qualified_request_cpu_jtag_debug_module,
      cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave => cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
      cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 => cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 => cpu_data_master_qualified_request_pio_bitcrusher_crush_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 => cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 => cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 => cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 => cpu_data_master_qualified_request_pio_bitcrusher_tone_s1,
      cpu_data_master_qualified_request_pio_compressor_bypass_s1 => cpu_data_master_qualified_request_pio_compressor_bypass_s1,
      cpu_data_master_qualified_request_pio_compressor_gain_s1 => cpu_data_master_qualified_request_pio_compressor_gain_s1,
      cpu_data_master_qualified_request_pio_compressor_treshold_s1 => cpu_data_master_qualified_request_pio_compressor_treshold_s1,
      cpu_data_master_qualified_request_pio_delay_bypass_s1 => cpu_data_master_qualified_request_pio_delay_bypass_s1,
      cpu_data_master_qualified_request_pio_delay_decay_s1 => cpu_data_master_qualified_request_pio_delay_decay_s1,
      cpu_data_master_qualified_request_pio_delay_length_s1 => cpu_data_master_qualified_request_pio_delay_length_s1,
      cpu_data_master_qualified_request_pio_master_volume_s1 => cpu_data_master_qualified_request_pio_master_volume_s1,
      cpu_data_master_qualified_request_pio_octaver_bypass_s1 => cpu_data_master_qualified_request_pio_octaver_bypass_s1,
      cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 => cpu_data_master_qualified_request_pio_octaver_dry_wet_s1,
      cpu_data_master_qualified_request_pio_output_power_left_s1 => cpu_data_master_qualified_request_pio_output_power_left_s1,
      cpu_data_master_qualified_request_pio_output_power_right_s1 => cpu_data_master_qualified_request_pio_output_power_right_s1,
      cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 => cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1,
      cpu_data_master_qualified_request_pio_overdrive_bypass_s1 => cpu_data_master_qualified_request_pio_overdrive_bypass_s1,
      cpu_data_master_qualified_request_pio_overdrive_gain_s1 => cpu_data_master_qualified_request_pio_overdrive_gain_s1,
      cpu_data_master_qualified_request_pio_overdrive_tone_s1 => cpu_data_master_qualified_request_pio_overdrive_tone_s1,
      cpu_data_master_qualified_request_pio_overdrive_volume_s1 => cpu_data_master_qualified_request_pio_overdrive_volume_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1,
      cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave,
      cpu_data_master_qualified_request_ps2_avalon_ps2_slave => cpu_data_master_qualified_request_ps2_avalon_ps2_slave,
      cpu_data_master_qualified_request_sdram_s1 => cpu_data_master_qualified_request_sdram_s1,
      cpu_data_master_qualified_request_sram_avalon_sram_slave => cpu_data_master_qualified_request_sram_avalon_sram_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_read_data_valid_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave => cpu_data_master_read_data_valid_analyzer_input_left_avalon_slave,
      cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave => cpu_data_master_read_data_valid_analyzer_input_right_avalon_slave,
      cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave,
      cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave => cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave => cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave,
      cpu_data_master_read_data_valid_cpu_jtag_debug_module => cpu_data_master_read_data_valid_cpu_jtag_debug_module,
      cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave => cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
      cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1,
      cpu_data_master_read_data_valid_pio_compressor_bypass_s1 => cpu_data_master_read_data_valid_pio_compressor_bypass_s1,
      cpu_data_master_read_data_valid_pio_compressor_gain_s1 => cpu_data_master_read_data_valid_pio_compressor_gain_s1,
      cpu_data_master_read_data_valid_pio_compressor_treshold_s1 => cpu_data_master_read_data_valid_pio_compressor_treshold_s1,
      cpu_data_master_read_data_valid_pio_delay_bypass_s1 => cpu_data_master_read_data_valid_pio_delay_bypass_s1,
      cpu_data_master_read_data_valid_pio_delay_decay_s1 => cpu_data_master_read_data_valid_pio_delay_decay_s1,
      cpu_data_master_read_data_valid_pio_delay_length_s1 => cpu_data_master_read_data_valid_pio_delay_length_s1,
      cpu_data_master_read_data_valid_pio_master_volume_s1 => cpu_data_master_read_data_valid_pio_master_volume_s1,
      cpu_data_master_read_data_valid_pio_octaver_bypass_s1 => cpu_data_master_read_data_valid_pio_octaver_bypass_s1,
      cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1 => cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1,
      cpu_data_master_read_data_valid_pio_output_power_left_s1 => cpu_data_master_read_data_valid_pio_output_power_left_s1,
      cpu_data_master_read_data_valid_pio_output_power_right_s1 => cpu_data_master_read_data_valid_pio_output_power_right_s1,
      cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1 => cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1,
      cpu_data_master_read_data_valid_pio_overdrive_bypass_s1 => cpu_data_master_read_data_valid_pio_overdrive_bypass_s1,
      cpu_data_master_read_data_valid_pio_overdrive_gain_s1 => cpu_data_master_read_data_valid_pio_overdrive_gain_s1,
      cpu_data_master_read_data_valid_pio_overdrive_tone_s1 => cpu_data_master_read_data_valid_pio_overdrive_tone_s1,
      cpu_data_master_read_data_valid_pio_overdrive_volume_s1 => cpu_data_master_read_data_valid_pio_overdrive_volume_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1,
      cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave,
      cpu_data_master_read_data_valid_ps2_avalon_ps2_slave => cpu_data_master_read_data_valid_ps2_avalon_ps2_slave,
      cpu_data_master_read_data_valid_sdram_s1 => cpu_data_master_read_data_valid_sdram_s1,
      cpu_data_master_read_data_valid_sdram_s1_shift_register => cpu_data_master_read_data_valid_sdram_s1_shift_register,
      cpu_data_master_read_data_valid_sram_avalon_sram_slave => cpu_data_master_read_data_valid_sram_avalon_sram_slave,
      cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data => cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data,
      cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control => cpu_data_master_requests_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control,
      cpu_data_master_requests_analyzer_input_left_avalon_slave => cpu_data_master_requests_analyzer_input_left_avalon_slave,
      cpu_data_master_requests_analyzer_input_right_avalon_slave => cpu_data_master_requests_analyzer_input_right_avalon_slave,
      cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave => cpu_data_master_requests_audio_and_video_config_0_avalon_on_board_config_slave,
      cpu_data_master_requests_character_buffer_avalon_char_buffer_slave => cpu_data_master_requests_character_buffer_avalon_char_buffer_slave,
      cpu_data_master_requests_character_buffer_avalon_char_control_slave => cpu_data_master_requests_character_buffer_avalon_char_control_slave,
      cpu_data_master_requests_cpu_jtag_debug_module => cpu_data_master_requests_cpu_jtag_debug_module,
      cpu_data_master_requests_jtag_uart_avalon_jtag_slave => cpu_data_master_requests_jtag_uart_avalon_jtag_slave,
      cpu_data_master_requests_pio_bitcrusher_bypass_s1 => cpu_data_master_requests_pio_bitcrusher_bypass_s1,
      cpu_data_master_requests_pio_bitcrusher_crush_s1 => cpu_data_master_requests_pio_bitcrusher_crush_s1,
      cpu_data_master_requests_pio_bitcrusher_downsample_s1 => cpu_data_master_requests_pio_bitcrusher_downsample_s1,
      cpu_data_master_requests_pio_bitcrusher_drywet_s1 => cpu_data_master_requests_pio_bitcrusher_drywet_s1,
      cpu_data_master_requests_pio_bitcrusher_flavor_s1 => cpu_data_master_requests_pio_bitcrusher_flavor_s1,
      cpu_data_master_requests_pio_bitcrusher_tone_s1 => cpu_data_master_requests_pio_bitcrusher_tone_s1,
      cpu_data_master_requests_pio_compressor_bypass_s1 => cpu_data_master_requests_pio_compressor_bypass_s1,
      cpu_data_master_requests_pio_compressor_gain_s1 => cpu_data_master_requests_pio_compressor_gain_s1,
      cpu_data_master_requests_pio_compressor_treshold_s1 => cpu_data_master_requests_pio_compressor_treshold_s1,
      cpu_data_master_requests_pio_delay_bypass_s1 => cpu_data_master_requests_pio_delay_bypass_s1,
      cpu_data_master_requests_pio_delay_decay_s1 => cpu_data_master_requests_pio_delay_decay_s1,
      cpu_data_master_requests_pio_delay_length_s1 => cpu_data_master_requests_pio_delay_length_s1,
      cpu_data_master_requests_pio_master_volume_s1 => cpu_data_master_requests_pio_master_volume_s1,
      cpu_data_master_requests_pio_octaver_bypass_s1 => cpu_data_master_requests_pio_octaver_bypass_s1,
      cpu_data_master_requests_pio_octaver_dry_wet_s1 => cpu_data_master_requests_pio_octaver_dry_wet_s1,
      cpu_data_master_requests_pio_output_power_left_s1 => cpu_data_master_requests_pio_output_power_left_s1,
      cpu_data_master_requests_pio_output_power_right_s1 => cpu_data_master_requests_pio_output_power_right_s1,
      cpu_data_master_requests_pio_overdrive_asymmetric_s1 => cpu_data_master_requests_pio_overdrive_asymmetric_s1,
      cpu_data_master_requests_pio_overdrive_bypass_s1 => cpu_data_master_requests_pio_overdrive_bypass_s1,
      cpu_data_master_requests_pio_overdrive_gain_s1 => cpu_data_master_requests_pio_overdrive_gain_s1,
      cpu_data_master_requests_pio_overdrive_tone_s1 => cpu_data_master_requests_pio_overdrive_tone_s1,
      cpu_data_master_requests_pio_overdrive_volume_s1 => cpu_data_master_requests_pio_overdrive_volume_s1,
      cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 => cpu_data_master_requests_pio_tremolo_stereo_bypass_s1,
      cpu_data_master_requests_pio_tremolo_stereo_depth_s1 => cpu_data_master_requests_pio_tremolo_stereo_depth_s1,
      cpu_data_master_requests_pio_tremolo_stereo_mode_s1 => cpu_data_master_requests_pio_tremolo_stereo_mode_s1,
      cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1,
      cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1,
      cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave,
      cpu_data_master_requests_ps2_avalon_ps2_slave => cpu_data_master_requests_ps2_avalon_ps2_slave,
      cpu_data_master_requests_sdram_s1 => cpu_data_master_requests_sdram_s1,
      cpu_data_master_requests_sram_avalon_sram_slave => cpu_data_master_requests_sram_avalon_sram_slave,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer => d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_end_xfer,
      d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer => d1_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_end_xfer,
      d1_analyzer_input_left_avalon_slave_end_xfer => d1_analyzer_input_left_avalon_slave_end_xfer,
      d1_analyzer_input_right_avalon_slave_end_xfer => d1_analyzer_input_right_avalon_slave_end_xfer,
      d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer => d1_audio_and_video_config_0_avalon_on_board_config_slave_end_xfer,
      d1_character_buffer_avalon_char_buffer_slave_end_xfer => d1_character_buffer_avalon_char_buffer_slave_end_xfer,
      d1_character_buffer_avalon_char_control_slave_end_xfer => d1_character_buffer_avalon_char_control_slave_end_xfer,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      d1_pio_bitcrusher_bypass_s1_end_xfer => d1_pio_bitcrusher_bypass_s1_end_xfer,
      d1_pio_bitcrusher_crush_s1_end_xfer => d1_pio_bitcrusher_crush_s1_end_xfer,
      d1_pio_bitcrusher_downsample_s1_end_xfer => d1_pio_bitcrusher_downsample_s1_end_xfer,
      d1_pio_bitcrusher_drywet_s1_end_xfer => d1_pio_bitcrusher_drywet_s1_end_xfer,
      d1_pio_bitcrusher_flavor_s1_end_xfer => d1_pio_bitcrusher_flavor_s1_end_xfer,
      d1_pio_bitcrusher_tone_s1_end_xfer => d1_pio_bitcrusher_tone_s1_end_xfer,
      d1_pio_compressor_bypass_s1_end_xfer => d1_pio_compressor_bypass_s1_end_xfer,
      d1_pio_compressor_gain_s1_end_xfer => d1_pio_compressor_gain_s1_end_xfer,
      d1_pio_compressor_treshold_s1_end_xfer => d1_pio_compressor_treshold_s1_end_xfer,
      d1_pio_delay_bypass_s1_end_xfer => d1_pio_delay_bypass_s1_end_xfer,
      d1_pio_delay_decay_s1_end_xfer => d1_pio_delay_decay_s1_end_xfer,
      d1_pio_delay_length_s1_end_xfer => d1_pio_delay_length_s1_end_xfer,
      d1_pio_master_volume_s1_end_xfer => d1_pio_master_volume_s1_end_xfer,
      d1_pio_octaver_bypass_s1_end_xfer => d1_pio_octaver_bypass_s1_end_xfer,
      d1_pio_octaver_dry_wet_s1_end_xfer => d1_pio_octaver_dry_wet_s1_end_xfer,
      d1_pio_output_power_left_s1_end_xfer => d1_pio_output_power_left_s1_end_xfer,
      d1_pio_output_power_right_s1_end_xfer => d1_pio_output_power_right_s1_end_xfer,
      d1_pio_overdrive_asymmetric_s1_end_xfer => d1_pio_overdrive_asymmetric_s1_end_xfer,
      d1_pio_overdrive_bypass_s1_end_xfer => d1_pio_overdrive_bypass_s1_end_xfer,
      d1_pio_overdrive_gain_s1_end_xfer => d1_pio_overdrive_gain_s1_end_xfer,
      d1_pio_overdrive_tone_s1_end_xfer => d1_pio_overdrive_tone_s1_end_xfer,
      d1_pio_overdrive_volume_s1_end_xfer => d1_pio_overdrive_volume_s1_end_xfer,
      d1_pio_tremolo_stereo_bypass_s1_end_xfer => d1_pio_tremolo_stereo_bypass_s1_end_xfer,
      d1_pio_tremolo_stereo_depth_s1_end_xfer => d1_pio_tremolo_stereo_depth_s1_end_xfer,
      d1_pio_tremolo_stereo_mode_s1_end_xfer => d1_pio_tremolo_stereo_mode_s1_end_xfer,
      d1_pio_tremolo_stereo_sweep_a_s1_end_xfer => d1_pio_tremolo_stereo_sweep_a_s1_end_xfer,
      d1_pio_tremolo_stereo_sweep_b_s1_end_xfer => d1_pio_tremolo_stereo_sweep_b_s1_end_xfer,
      d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer => d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer,
      d1_ps2_avalon_ps2_slave_end_xfer => d1_ps2_avalon_ps2_slave_end_xfer,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      d1_sram_avalon_sram_slave_end_xfer => d1_sram_avalon_sram_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      pio_bitcrusher_bypass_s1_readdata_from_sa => pio_bitcrusher_bypass_s1_readdata_from_sa,
      pio_bitcrusher_crush_s1_readdata_from_sa => pio_bitcrusher_crush_s1_readdata_from_sa,
      pio_bitcrusher_downsample_s1_readdata_from_sa => pio_bitcrusher_downsample_s1_readdata_from_sa,
      pio_bitcrusher_drywet_s1_readdata_from_sa => pio_bitcrusher_drywet_s1_readdata_from_sa,
      pio_bitcrusher_flavor_s1_readdata_from_sa => pio_bitcrusher_flavor_s1_readdata_from_sa,
      pio_bitcrusher_tone_s1_readdata_from_sa => pio_bitcrusher_tone_s1_readdata_from_sa,
      pio_compressor_bypass_s1_readdata_from_sa => pio_compressor_bypass_s1_readdata_from_sa,
      pio_compressor_gain_s1_readdata_from_sa => pio_compressor_gain_s1_readdata_from_sa,
      pio_compressor_treshold_s1_readdata_from_sa => pio_compressor_treshold_s1_readdata_from_sa,
      pio_delay_bypass_s1_readdata_from_sa => pio_delay_bypass_s1_readdata_from_sa,
      pio_delay_decay_s1_readdata_from_sa => pio_delay_decay_s1_readdata_from_sa,
      pio_delay_length_s1_readdata_from_sa => pio_delay_length_s1_readdata_from_sa,
      pio_master_volume_s1_readdata_from_sa => pio_master_volume_s1_readdata_from_sa,
      pio_octaver_bypass_s1_readdata_from_sa => pio_octaver_bypass_s1_readdata_from_sa,
      pio_octaver_dry_wet_s1_readdata_from_sa => pio_octaver_dry_wet_s1_readdata_from_sa,
      pio_output_power_left_s1_readdata_from_sa => pio_output_power_left_s1_readdata_from_sa,
      pio_output_power_right_s1_readdata_from_sa => pio_output_power_right_s1_readdata_from_sa,
      pio_overdrive_asymmetric_s1_readdata_from_sa => pio_overdrive_asymmetric_s1_readdata_from_sa,
      pio_overdrive_bypass_s1_readdata_from_sa => pio_overdrive_bypass_s1_readdata_from_sa,
      pio_overdrive_gain_s1_readdata_from_sa => pio_overdrive_gain_s1_readdata_from_sa,
      pio_overdrive_tone_s1_readdata_from_sa => pio_overdrive_tone_s1_readdata_from_sa,
      pio_overdrive_volume_s1_readdata_from_sa => pio_overdrive_volume_s1_readdata_from_sa,
      pio_tremolo_stereo_bypass_s1_readdata_from_sa => pio_tremolo_stereo_bypass_s1_readdata_from_sa,
      pio_tremolo_stereo_depth_s1_readdata_from_sa => pio_tremolo_stereo_depth_s1_readdata_from_sa,
      pio_tremolo_stereo_mode_s1_readdata_from_sa => pio_tremolo_stereo_mode_s1_readdata_from_sa,
      pio_tremolo_stereo_sweep_a_s1_readdata_from_sa => pio_tremolo_stereo_sweep_a_s1_readdata_from_sa,
      pio_tremolo_stereo_sweep_b_s1_readdata_from_sa => pio_tremolo_stereo_sweep_b_s1_readdata_from_sa,
      pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa => pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa,
      ps2_avalon_ps2_slave_irq_from_sa => ps2_avalon_ps2_slave_irq_from_sa,
      ps2_avalon_ps2_slave_readdata_from_sa => ps2_avalon_ps2_slave_readdata_from_sa,
      ps2_avalon_ps2_slave_waitrequest_from_sa => ps2_avalon_ps2_slave_waitrequest_from_sa,
      registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave => registered_cpu_data_master_read_data_valid_audio_and_video_config_0_avalon_on_board_config_slave,
      registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave => registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_buffer_slave,
      registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave => registered_cpu_data_master_read_data_valid_character_buffer_avalon_char_control_slave,
      registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave => registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave,
      registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave => registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave,
      registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave => registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave,
      reset_n => clk_0_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa,
      sram_avalon_sram_slave_readdata_from_sa => sram_avalon_sram_slave_readdata_from_sa
    );


  --the_cpu_instruction_master, which is an e_instance
  the_cpu_instruction_master : cpu_instruction_master_arbitrator
    port map(
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_dbs_address => cpu_instruction_master_dbs_address,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_readdata => cpu_instruction_master_readdata,
      cpu_instruction_master_readdatavalid => cpu_instruction_master_readdatavalid,
      cpu_instruction_master_waitrequest => cpu_instruction_master_waitrequest,
      clk => clk_0,
      cpu_instruction_master_address => cpu_instruction_master_address,
      cpu_instruction_master_granted_cpu_jtag_debug_module => cpu_instruction_master_granted_cpu_jtag_debug_module,
      cpu_instruction_master_granted_sram_avalon_sram_slave => cpu_instruction_master_granted_sram_avalon_sram_slave,
      cpu_instruction_master_qualified_request_cpu_jtag_debug_module => cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
      cpu_instruction_master_qualified_request_sram_avalon_sram_slave => cpu_instruction_master_qualified_request_sram_avalon_sram_slave,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_cpu_jtag_debug_module => cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
      cpu_instruction_master_read_data_valid_sram_avalon_sram_slave => cpu_instruction_master_read_data_valid_sram_avalon_sram_slave,
      cpu_instruction_master_requests_cpu_jtag_debug_module => cpu_instruction_master_requests_cpu_jtag_debug_module,
      cpu_instruction_master_requests_sram_avalon_sram_slave => cpu_instruction_master_requests_sram_avalon_sram_slave,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      d1_sram_avalon_sram_slave_end_xfer => d1_sram_avalon_sram_slave_end_xfer,
      reset_n => clk_0_reset_n,
      sram_avalon_sram_slave_readdata_from_sa => sram_avalon_sram_slave_readdata_from_sa
    );


  --the_cpu, which is an e_ptf_instance
  the_cpu : cpu
    port map(
      A_ci_multi_a => cpu_custom_instruction_master_multi_a,
      A_ci_multi_b => cpu_custom_instruction_master_multi_b,
      A_ci_multi_c => cpu_custom_instruction_master_multi_c,
      A_ci_multi_clk_en => cpu_custom_instruction_master_multi_clk_en,
      A_ci_multi_dataa => cpu_custom_instruction_master_multi_dataa,
      A_ci_multi_datab => cpu_custom_instruction_master_multi_datab,
      A_ci_multi_estatus => cpu_custom_instruction_master_multi_estatus,
      A_ci_multi_ipending => cpu_custom_instruction_master_multi_ipending,
      A_ci_multi_n => cpu_custom_instruction_master_multi_n,
      A_ci_multi_readra => cpu_custom_instruction_master_multi_readra,
      A_ci_multi_readrb => cpu_custom_instruction_master_multi_readrb,
      A_ci_multi_start => cpu_custom_instruction_master_multi_start,
      A_ci_multi_status => cpu_custom_instruction_master_multi_status,
      A_ci_multi_writerc => cpu_custom_instruction_master_multi_writerc,
      d_address => cpu_data_master_address,
      d_byteenable => cpu_data_master_byteenable,
      d_read => cpu_data_master_read,
      d_write => cpu_data_master_write,
      d_writedata => cpu_data_master_writedata,
      i_address => cpu_instruction_master_address,
      i_read => cpu_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,
      jtag_debug_module_readdata => cpu_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => cpu_jtag_debug_module_resetrequest,
      A_ci_multi_done => cpu_custom_instruction_master_multi_done,
      A_ci_multi_result => cpu_custom_instruction_master_multi_result,
      clk => clk_0,
      d_irq => cpu_data_master_irq,
      d_readdata => cpu_data_master_readdata,
      d_waitrequest => cpu_data_master_waitrequest,
      i_readdata => cpu_instruction_master_readdata,
      i_readdatavalid => cpu_instruction_master_readdatavalid,
      i_waitrequest => cpu_instruction_master_waitrequest,
      jtag_debug_module_address => cpu_jtag_debug_module_address,
      jtag_debug_module_begintransfer => cpu_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => cpu_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => cpu_jtag_debug_module_debugaccess,
      jtag_debug_module_select => cpu_jtag_debug_module_chipselect,
      jtag_debug_module_write => cpu_jtag_debug_module_write,
      jtag_debug_module_writedata => cpu_jtag_debug_module_writedata,
      reset_n => cpu_custom_instruction_master_reset_n
    );


  --the_cpu_fpoint_s1, which is an e_instance
  the_cpu_fpoint_s1 : cpu_fpoint_s1_arbitrator
    port map(
      cpu_fpoint_s1_clk_en => cpu_fpoint_s1_clk_en,
      cpu_fpoint_s1_dataa => cpu_fpoint_s1_dataa,
      cpu_fpoint_s1_datab => cpu_fpoint_s1_datab,
      cpu_fpoint_s1_done_from_sa => cpu_fpoint_s1_done_from_sa,
      cpu_fpoint_s1_n => cpu_fpoint_s1_n,
      cpu_fpoint_s1_reset => cpu_fpoint_s1_reset,
      cpu_fpoint_s1_result_from_sa => cpu_fpoint_s1_result_from_sa,
      cpu_fpoint_s1_start => cpu_fpoint_s1_start,
      clk => clk_0,
      cpu_custom_instruction_master_multi_clk_en => cpu_custom_instruction_master_multi_clk_en,
      cpu_custom_instruction_master_multi_dataa => cpu_custom_instruction_master_multi_dataa,
      cpu_custom_instruction_master_multi_datab => cpu_custom_instruction_master_multi_datab,
      cpu_custom_instruction_master_multi_n => cpu_custom_instruction_master_multi_n,
      cpu_custom_instruction_master_start_cpu_fpoint_s1 => cpu_custom_instruction_master_start_cpu_fpoint_s1,
      cpu_fpoint_s1_done => cpu_fpoint_s1_done,
      cpu_fpoint_s1_result => cpu_fpoint_s1_result,
      cpu_fpoint_s1_select => cpu_fpoint_s1_select,
      reset_n => clk_0_reset_n
    );


  --the_cpu_fpoint, which is an e_ptf_instance
  the_cpu_fpoint : cpu_fpoint
    port map(
      done => cpu_fpoint_s1_done,
      result => cpu_fpoint_s1_result,
      clk => clk_0,
      clk_en => cpu_fpoint_s1_clk_en,
      dataa => cpu_fpoint_s1_dataa,
      datab => cpu_fpoint_s1_datab,
      n => cpu_fpoint_s1_n,
      reset => cpu_fpoint_s1_reset,
      start => cpu_fpoint_s1_start
    );


  --the_jtag_uart_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_avalon_jtag_slave : jtag_uart_avalon_jtag_slave_arbitrator
    port map(
      cpu_data_master_granted_jtag_uart_avalon_jtag_slave => cpu_data_master_granted_jtag_uart_avalon_jtag_slave,
      cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave => cpu_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
      cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave => cpu_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
      cpu_data_master_requests_jtag_uart_avalon_jtag_slave => cpu_data_master_requests_jtag_uart_avalon_jtag_slave,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_address => jtag_uart_avalon_jtag_slave_address,
      jtag_uart_avalon_jtag_slave_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      jtag_uart_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_read_n => jtag_uart_avalon_jtag_slave_read_n,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_avalon_jtag_slave_reset_n => jtag_uart_avalon_jtag_slave_reset_n,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_avalon_jtag_slave_write_n => jtag_uart_avalon_jtag_slave_write_n,
      jtag_uart_avalon_jtag_slave_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      jtag_uart_avalon_jtag_slave_dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      jtag_uart_avalon_jtag_slave_irq => jtag_uart_avalon_jtag_slave_irq,
      jtag_uart_avalon_jtag_slave_readdata => jtag_uart_avalon_jtag_slave_readdata,
      jtag_uart_avalon_jtag_slave_readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      jtag_uart_avalon_jtag_slave_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      reset_n => clk_0_reset_n
    );


  --the_jtag_uart, which is an e_ptf_instance
  the_jtag_uart : jtag_uart
    port map(
      av_irq => jtag_uart_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => clk_0,
      rst_n => jtag_uart_avalon_jtag_slave_reset_n
    );


  --the_membuffer_0_avalon_master, which is an e_instance
  the_membuffer_0_avalon_master : membuffer_0_avalon_master_arbitrator
    port map(
      membuffer_0_avalon_master_address_to_slave => membuffer_0_avalon_master_address_to_slave,
      membuffer_0_avalon_master_readdata => membuffer_0_avalon_master_readdata,
      membuffer_0_avalon_master_reset_n => membuffer_0_avalon_master_reset_n,
      membuffer_0_avalon_master_waitrequest => membuffer_0_avalon_master_waitrequest,
      membuffer_0_dbs_address => membuffer_0_dbs_address,
      membuffer_0_dbs_write_16 => membuffer_0_dbs_write_16,
      clk => clk_0,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      membuffer_0_avalon_master_address => membuffer_0_avalon_master_address,
      membuffer_0_avalon_master_read => membuffer_0_avalon_master_read,
      membuffer_0_avalon_master_write => membuffer_0_avalon_master_write,
      membuffer_0_avalon_master_writedata => membuffer_0_avalon_master_writedata,
      membuffer_0_byteenable_sdram_s1 => membuffer_0_byteenable_sdram_s1,
      membuffer_0_granted_sdram_s1 => membuffer_0_granted_sdram_s1,
      membuffer_0_qualified_request_sdram_s1 => membuffer_0_qualified_request_sdram_s1,
      membuffer_0_read_data_valid_sdram_s1 => membuffer_0_read_data_valid_sdram_s1,
      membuffer_0_read_data_valid_sdram_s1_shift_register => membuffer_0_read_data_valid_sdram_s1_shift_register,
      membuffer_0_requests_sdram_s1 => membuffer_0_requests_sdram_s1,
      reset_n => clk_0_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_membuffer_0, which is an e_ptf_instance
  the_membuffer_0 : membuffer_0
    port map(
      address => membuffer_0_avalon_master_address,
      read => membuffer_0_avalon_master_read,
      sample_left_out => internal_sample_left_out_from_the_membuffer_0,
      sample_right_out => internal_sample_right_out_from_the_membuffer_0,
      write => membuffer_0_avalon_master_write,
      writedata => membuffer_0_avalon_master_writedata,
      clk => clk_0,
      delay_time => delay_time_to_the_membuffer_0,
      readdata => membuffer_0_avalon_master_readdata,
      reset => membuffer_0_avalon_master_reset_n,
      sample_clk => sample_clk_to_the_membuffer_0,
      sample_left_in => sample_left_in_to_the_membuffer_0,
      sample_right_in => sample_right_in_to_the_membuffer_0,
      waitrequest => membuffer_0_avalon_master_waitrequest
    );


  --the_pio_bitcrusher_bypass_s1, which is an e_instance
  the_pio_bitcrusher_bypass_s1 : pio_bitcrusher_bypass_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_bitcrusher_bypass_s1 => cpu_data_master_granted_pio_bitcrusher_bypass_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1 => cpu_data_master_qualified_request_pio_bitcrusher_bypass_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_bypass_s1,
      cpu_data_master_requests_pio_bitcrusher_bypass_s1 => cpu_data_master_requests_pio_bitcrusher_bypass_s1,
      d1_pio_bitcrusher_bypass_s1_end_xfer => d1_pio_bitcrusher_bypass_s1_end_xfer,
      pio_bitcrusher_bypass_s1_address => pio_bitcrusher_bypass_s1_address,
      pio_bitcrusher_bypass_s1_chipselect => pio_bitcrusher_bypass_s1_chipselect,
      pio_bitcrusher_bypass_s1_readdata_from_sa => pio_bitcrusher_bypass_s1_readdata_from_sa,
      pio_bitcrusher_bypass_s1_reset_n => pio_bitcrusher_bypass_s1_reset_n,
      pio_bitcrusher_bypass_s1_write_n => pio_bitcrusher_bypass_s1_write_n,
      pio_bitcrusher_bypass_s1_writedata => pio_bitcrusher_bypass_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_bitcrusher_bypass_s1_readdata => pio_bitcrusher_bypass_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_bitcrusher_bypass, which is an e_ptf_instance
  the_pio_bitcrusher_bypass : pio_bitcrusher_bypass
    port map(
      out_port => internal_out_port_from_the_pio_bitcrusher_bypass,
      readdata => pio_bitcrusher_bypass_s1_readdata,
      address => pio_bitcrusher_bypass_s1_address,
      chipselect => pio_bitcrusher_bypass_s1_chipselect,
      clk => clk_0,
      reset_n => pio_bitcrusher_bypass_s1_reset_n,
      write_n => pio_bitcrusher_bypass_s1_write_n,
      writedata => pio_bitcrusher_bypass_s1_writedata
    );


  --the_pio_bitcrusher_crush_s1, which is an e_instance
  the_pio_bitcrusher_crush_s1 : pio_bitcrusher_crush_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_bitcrusher_crush_s1 => cpu_data_master_granted_pio_bitcrusher_crush_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_crush_s1 => cpu_data_master_qualified_request_pio_bitcrusher_crush_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_crush_s1,
      cpu_data_master_requests_pio_bitcrusher_crush_s1 => cpu_data_master_requests_pio_bitcrusher_crush_s1,
      d1_pio_bitcrusher_crush_s1_end_xfer => d1_pio_bitcrusher_crush_s1_end_xfer,
      pio_bitcrusher_crush_s1_address => pio_bitcrusher_crush_s1_address,
      pio_bitcrusher_crush_s1_chipselect => pio_bitcrusher_crush_s1_chipselect,
      pio_bitcrusher_crush_s1_readdata_from_sa => pio_bitcrusher_crush_s1_readdata_from_sa,
      pio_bitcrusher_crush_s1_reset_n => pio_bitcrusher_crush_s1_reset_n,
      pio_bitcrusher_crush_s1_write_n => pio_bitcrusher_crush_s1_write_n,
      pio_bitcrusher_crush_s1_writedata => pio_bitcrusher_crush_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_bitcrusher_crush_s1_readdata => pio_bitcrusher_crush_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_bitcrusher_crush, which is an e_ptf_instance
  the_pio_bitcrusher_crush : pio_bitcrusher_crush
    port map(
      out_port => internal_out_port_from_the_pio_bitcrusher_crush,
      readdata => pio_bitcrusher_crush_s1_readdata,
      address => pio_bitcrusher_crush_s1_address,
      chipselect => pio_bitcrusher_crush_s1_chipselect,
      clk => clk_0,
      reset_n => pio_bitcrusher_crush_s1_reset_n,
      write_n => pio_bitcrusher_crush_s1_write_n,
      writedata => pio_bitcrusher_crush_s1_writedata
    );


  --the_pio_bitcrusher_downsample_s1, which is an e_instance
  the_pio_bitcrusher_downsample_s1 : pio_bitcrusher_downsample_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_bitcrusher_downsample_s1 => cpu_data_master_granted_pio_bitcrusher_downsample_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1 => cpu_data_master_qualified_request_pio_bitcrusher_downsample_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_downsample_s1,
      cpu_data_master_requests_pio_bitcrusher_downsample_s1 => cpu_data_master_requests_pio_bitcrusher_downsample_s1,
      d1_pio_bitcrusher_downsample_s1_end_xfer => d1_pio_bitcrusher_downsample_s1_end_xfer,
      pio_bitcrusher_downsample_s1_address => pio_bitcrusher_downsample_s1_address,
      pio_bitcrusher_downsample_s1_chipselect => pio_bitcrusher_downsample_s1_chipselect,
      pio_bitcrusher_downsample_s1_readdata_from_sa => pio_bitcrusher_downsample_s1_readdata_from_sa,
      pio_bitcrusher_downsample_s1_reset_n => pio_bitcrusher_downsample_s1_reset_n,
      pio_bitcrusher_downsample_s1_write_n => pio_bitcrusher_downsample_s1_write_n,
      pio_bitcrusher_downsample_s1_writedata => pio_bitcrusher_downsample_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_bitcrusher_downsample_s1_readdata => pio_bitcrusher_downsample_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_bitcrusher_downsample, which is an e_ptf_instance
  the_pio_bitcrusher_downsample : pio_bitcrusher_downsample
    port map(
      out_port => internal_out_port_from_the_pio_bitcrusher_downsample,
      readdata => pio_bitcrusher_downsample_s1_readdata,
      address => pio_bitcrusher_downsample_s1_address,
      chipselect => pio_bitcrusher_downsample_s1_chipselect,
      clk => clk_0,
      reset_n => pio_bitcrusher_downsample_s1_reset_n,
      write_n => pio_bitcrusher_downsample_s1_write_n,
      writedata => pio_bitcrusher_downsample_s1_writedata
    );


  --the_pio_bitcrusher_drywet_s1, which is an e_instance
  the_pio_bitcrusher_drywet_s1 : pio_bitcrusher_drywet_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_bitcrusher_drywet_s1 => cpu_data_master_granted_pio_bitcrusher_drywet_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1 => cpu_data_master_qualified_request_pio_bitcrusher_drywet_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_drywet_s1,
      cpu_data_master_requests_pio_bitcrusher_drywet_s1 => cpu_data_master_requests_pio_bitcrusher_drywet_s1,
      d1_pio_bitcrusher_drywet_s1_end_xfer => d1_pio_bitcrusher_drywet_s1_end_xfer,
      pio_bitcrusher_drywet_s1_address => pio_bitcrusher_drywet_s1_address,
      pio_bitcrusher_drywet_s1_chipselect => pio_bitcrusher_drywet_s1_chipselect,
      pio_bitcrusher_drywet_s1_readdata_from_sa => pio_bitcrusher_drywet_s1_readdata_from_sa,
      pio_bitcrusher_drywet_s1_reset_n => pio_bitcrusher_drywet_s1_reset_n,
      pio_bitcrusher_drywet_s1_write_n => pio_bitcrusher_drywet_s1_write_n,
      pio_bitcrusher_drywet_s1_writedata => pio_bitcrusher_drywet_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_bitcrusher_drywet_s1_readdata => pio_bitcrusher_drywet_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_bitcrusher_drywet, which is an e_ptf_instance
  the_pio_bitcrusher_drywet : pio_bitcrusher_drywet
    port map(
      out_port => internal_out_port_from_the_pio_bitcrusher_drywet,
      readdata => pio_bitcrusher_drywet_s1_readdata,
      address => pio_bitcrusher_drywet_s1_address,
      chipselect => pio_bitcrusher_drywet_s1_chipselect,
      clk => clk_0,
      reset_n => pio_bitcrusher_drywet_s1_reset_n,
      write_n => pio_bitcrusher_drywet_s1_write_n,
      writedata => pio_bitcrusher_drywet_s1_writedata
    );


  --the_pio_bitcrusher_flavor_s1, which is an e_instance
  the_pio_bitcrusher_flavor_s1 : pio_bitcrusher_flavor_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_bitcrusher_flavor_s1 => cpu_data_master_granted_pio_bitcrusher_flavor_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1 => cpu_data_master_qualified_request_pio_bitcrusher_flavor_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_flavor_s1,
      cpu_data_master_requests_pio_bitcrusher_flavor_s1 => cpu_data_master_requests_pio_bitcrusher_flavor_s1,
      d1_pio_bitcrusher_flavor_s1_end_xfer => d1_pio_bitcrusher_flavor_s1_end_xfer,
      pio_bitcrusher_flavor_s1_address => pio_bitcrusher_flavor_s1_address,
      pio_bitcrusher_flavor_s1_chipselect => pio_bitcrusher_flavor_s1_chipselect,
      pio_bitcrusher_flavor_s1_readdata_from_sa => pio_bitcrusher_flavor_s1_readdata_from_sa,
      pio_bitcrusher_flavor_s1_reset_n => pio_bitcrusher_flavor_s1_reset_n,
      pio_bitcrusher_flavor_s1_write_n => pio_bitcrusher_flavor_s1_write_n,
      pio_bitcrusher_flavor_s1_writedata => pio_bitcrusher_flavor_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_bitcrusher_flavor_s1_readdata => pio_bitcrusher_flavor_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_bitcrusher_flavor, which is an e_ptf_instance
  the_pio_bitcrusher_flavor : pio_bitcrusher_flavor
    port map(
      out_port => internal_out_port_from_the_pio_bitcrusher_flavor,
      readdata => pio_bitcrusher_flavor_s1_readdata,
      address => pio_bitcrusher_flavor_s1_address,
      chipselect => pio_bitcrusher_flavor_s1_chipselect,
      clk => clk_0,
      reset_n => pio_bitcrusher_flavor_s1_reset_n,
      write_n => pio_bitcrusher_flavor_s1_write_n,
      writedata => pio_bitcrusher_flavor_s1_writedata
    );


  --the_pio_bitcrusher_tone_s1, which is an e_instance
  the_pio_bitcrusher_tone_s1 : pio_bitcrusher_tone_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_bitcrusher_tone_s1 => cpu_data_master_granted_pio_bitcrusher_tone_s1,
      cpu_data_master_qualified_request_pio_bitcrusher_tone_s1 => cpu_data_master_qualified_request_pio_bitcrusher_tone_s1,
      cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1 => cpu_data_master_read_data_valid_pio_bitcrusher_tone_s1,
      cpu_data_master_requests_pio_bitcrusher_tone_s1 => cpu_data_master_requests_pio_bitcrusher_tone_s1,
      d1_pio_bitcrusher_tone_s1_end_xfer => d1_pio_bitcrusher_tone_s1_end_xfer,
      pio_bitcrusher_tone_s1_address => pio_bitcrusher_tone_s1_address,
      pio_bitcrusher_tone_s1_chipselect => pio_bitcrusher_tone_s1_chipselect,
      pio_bitcrusher_tone_s1_readdata_from_sa => pio_bitcrusher_tone_s1_readdata_from_sa,
      pio_bitcrusher_tone_s1_reset_n => pio_bitcrusher_tone_s1_reset_n,
      pio_bitcrusher_tone_s1_write_n => pio_bitcrusher_tone_s1_write_n,
      pio_bitcrusher_tone_s1_writedata => pio_bitcrusher_tone_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_bitcrusher_tone_s1_readdata => pio_bitcrusher_tone_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_bitcrusher_tone, which is an e_ptf_instance
  the_pio_bitcrusher_tone : pio_bitcrusher_tone
    port map(
      out_port => internal_out_port_from_the_pio_bitcrusher_tone,
      readdata => pio_bitcrusher_tone_s1_readdata,
      address => pio_bitcrusher_tone_s1_address,
      chipselect => pio_bitcrusher_tone_s1_chipselect,
      clk => clk_0,
      reset_n => pio_bitcrusher_tone_s1_reset_n,
      write_n => pio_bitcrusher_tone_s1_write_n,
      writedata => pio_bitcrusher_tone_s1_writedata
    );


  --the_pio_compressor_bypass_s1, which is an e_instance
  the_pio_compressor_bypass_s1 : pio_compressor_bypass_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_compressor_bypass_s1 => cpu_data_master_granted_pio_compressor_bypass_s1,
      cpu_data_master_qualified_request_pio_compressor_bypass_s1 => cpu_data_master_qualified_request_pio_compressor_bypass_s1,
      cpu_data_master_read_data_valid_pio_compressor_bypass_s1 => cpu_data_master_read_data_valid_pio_compressor_bypass_s1,
      cpu_data_master_requests_pio_compressor_bypass_s1 => cpu_data_master_requests_pio_compressor_bypass_s1,
      d1_pio_compressor_bypass_s1_end_xfer => d1_pio_compressor_bypass_s1_end_xfer,
      pio_compressor_bypass_s1_address => pio_compressor_bypass_s1_address,
      pio_compressor_bypass_s1_chipselect => pio_compressor_bypass_s1_chipselect,
      pio_compressor_bypass_s1_readdata_from_sa => pio_compressor_bypass_s1_readdata_from_sa,
      pio_compressor_bypass_s1_reset_n => pio_compressor_bypass_s1_reset_n,
      pio_compressor_bypass_s1_write_n => pio_compressor_bypass_s1_write_n,
      pio_compressor_bypass_s1_writedata => pio_compressor_bypass_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_compressor_bypass_s1_readdata => pio_compressor_bypass_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_compressor_bypass, which is an e_ptf_instance
  the_pio_compressor_bypass : pio_compressor_bypass
    port map(
      out_port => internal_out_port_from_the_pio_compressor_bypass,
      readdata => pio_compressor_bypass_s1_readdata,
      address => pio_compressor_bypass_s1_address,
      chipselect => pio_compressor_bypass_s1_chipselect,
      clk => clk_0,
      reset_n => pio_compressor_bypass_s1_reset_n,
      write_n => pio_compressor_bypass_s1_write_n,
      writedata => pio_compressor_bypass_s1_writedata
    );


  --the_pio_compressor_gain_s1, which is an e_instance
  the_pio_compressor_gain_s1 : pio_compressor_gain_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_compressor_gain_s1 => cpu_data_master_granted_pio_compressor_gain_s1,
      cpu_data_master_qualified_request_pio_compressor_gain_s1 => cpu_data_master_qualified_request_pio_compressor_gain_s1,
      cpu_data_master_read_data_valid_pio_compressor_gain_s1 => cpu_data_master_read_data_valid_pio_compressor_gain_s1,
      cpu_data_master_requests_pio_compressor_gain_s1 => cpu_data_master_requests_pio_compressor_gain_s1,
      d1_pio_compressor_gain_s1_end_xfer => d1_pio_compressor_gain_s1_end_xfer,
      pio_compressor_gain_s1_address => pio_compressor_gain_s1_address,
      pio_compressor_gain_s1_chipselect => pio_compressor_gain_s1_chipselect,
      pio_compressor_gain_s1_readdata_from_sa => pio_compressor_gain_s1_readdata_from_sa,
      pio_compressor_gain_s1_reset_n => pio_compressor_gain_s1_reset_n,
      pio_compressor_gain_s1_write_n => pio_compressor_gain_s1_write_n,
      pio_compressor_gain_s1_writedata => pio_compressor_gain_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_compressor_gain_s1_readdata => pio_compressor_gain_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_compressor_gain, which is an e_ptf_instance
  the_pio_compressor_gain : pio_compressor_gain
    port map(
      out_port => internal_out_port_from_the_pio_compressor_gain,
      readdata => pio_compressor_gain_s1_readdata,
      address => pio_compressor_gain_s1_address,
      chipselect => pio_compressor_gain_s1_chipselect,
      clk => clk_0,
      reset_n => pio_compressor_gain_s1_reset_n,
      write_n => pio_compressor_gain_s1_write_n,
      writedata => pio_compressor_gain_s1_writedata
    );


  --the_pio_compressor_treshold_s1, which is an e_instance
  the_pio_compressor_treshold_s1 : pio_compressor_treshold_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_compressor_treshold_s1 => cpu_data_master_granted_pio_compressor_treshold_s1,
      cpu_data_master_qualified_request_pio_compressor_treshold_s1 => cpu_data_master_qualified_request_pio_compressor_treshold_s1,
      cpu_data_master_read_data_valid_pio_compressor_treshold_s1 => cpu_data_master_read_data_valid_pio_compressor_treshold_s1,
      cpu_data_master_requests_pio_compressor_treshold_s1 => cpu_data_master_requests_pio_compressor_treshold_s1,
      d1_pio_compressor_treshold_s1_end_xfer => d1_pio_compressor_treshold_s1_end_xfer,
      pio_compressor_treshold_s1_address => pio_compressor_treshold_s1_address,
      pio_compressor_treshold_s1_chipselect => pio_compressor_treshold_s1_chipselect,
      pio_compressor_treshold_s1_readdata_from_sa => pio_compressor_treshold_s1_readdata_from_sa,
      pio_compressor_treshold_s1_reset_n => pio_compressor_treshold_s1_reset_n,
      pio_compressor_treshold_s1_write_n => pio_compressor_treshold_s1_write_n,
      pio_compressor_treshold_s1_writedata => pio_compressor_treshold_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_compressor_treshold_s1_readdata => pio_compressor_treshold_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_compressor_treshold, which is an e_ptf_instance
  the_pio_compressor_treshold : pio_compressor_treshold
    port map(
      out_port => internal_out_port_from_the_pio_compressor_treshold,
      readdata => pio_compressor_treshold_s1_readdata,
      address => pio_compressor_treshold_s1_address,
      chipselect => pio_compressor_treshold_s1_chipselect,
      clk => clk_0,
      reset_n => pio_compressor_treshold_s1_reset_n,
      write_n => pio_compressor_treshold_s1_write_n,
      writedata => pio_compressor_treshold_s1_writedata
    );


  --the_pio_delay_bypass_s1, which is an e_instance
  the_pio_delay_bypass_s1 : pio_delay_bypass_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_delay_bypass_s1 => cpu_data_master_granted_pio_delay_bypass_s1,
      cpu_data_master_qualified_request_pio_delay_bypass_s1 => cpu_data_master_qualified_request_pio_delay_bypass_s1,
      cpu_data_master_read_data_valid_pio_delay_bypass_s1 => cpu_data_master_read_data_valid_pio_delay_bypass_s1,
      cpu_data_master_requests_pio_delay_bypass_s1 => cpu_data_master_requests_pio_delay_bypass_s1,
      d1_pio_delay_bypass_s1_end_xfer => d1_pio_delay_bypass_s1_end_xfer,
      pio_delay_bypass_s1_address => pio_delay_bypass_s1_address,
      pio_delay_bypass_s1_chipselect => pio_delay_bypass_s1_chipselect,
      pio_delay_bypass_s1_readdata_from_sa => pio_delay_bypass_s1_readdata_from_sa,
      pio_delay_bypass_s1_reset_n => pio_delay_bypass_s1_reset_n,
      pio_delay_bypass_s1_write_n => pio_delay_bypass_s1_write_n,
      pio_delay_bypass_s1_writedata => pio_delay_bypass_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_delay_bypass_s1_readdata => pio_delay_bypass_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_delay_bypass, which is an e_ptf_instance
  the_pio_delay_bypass : pio_delay_bypass
    port map(
      out_port => internal_out_port_from_the_pio_delay_bypass,
      readdata => pio_delay_bypass_s1_readdata,
      address => pio_delay_bypass_s1_address,
      chipselect => pio_delay_bypass_s1_chipselect,
      clk => clk_0,
      reset_n => pio_delay_bypass_s1_reset_n,
      write_n => pio_delay_bypass_s1_write_n,
      writedata => pio_delay_bypass_s1_writedata
    );


  --the_pio_delay_decay_s1, which is an e_instance
  the_pio_delay_decay_s1 : pio_delay_decay_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_delay_decay_s1 => cpu_data_master_granted_pio_delay_decay_s1,
      cpu_data_master_qualified_request_pio_delay_decay_s1 => cpu_data_master_qualified_request_pio_delay_decay_s1,
      cpu_data_master_read_data_valid_pio_delay_decay_s1 => cpu_data_master_read_data_valid_pio_delay_decay_s1,
      cpu_data_master_requests_pio_delay_decay_s1 => cpu_data_master_requests_pio_delay_decay_s1,
      d1_pio_delay_decay_s1_end_xfer => d1_pio_delay_decay_s1_end_xfer,
      pio_delay_decay_s1_address => pio_delay_decay_s1_address,
      pio_delay_decay_s1_chipselect => pio_delay_decay_s1_chipselect,
      pio_delay_decay_s1_readdata_from_sa => pio_delay_decay_s1_readdata_from_sa,
      pio_delay_decay_s1_reset_n => pio_delay_decay_s1_reset_n,
      pio_delay_decay_s1_write_n => pio_delay_decay_s1_write_n,
      pio_delay_decay_s1_writedata => pio_delay_decay_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_delay_decay_s1_readdata => pio_delay_decay_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_delay_decay, which is an e_ptf_instance
  the_pio_delay_decay : pio_delay_decay
    port map(
      out_port => internal_out_port_from_the_pio_delay_decay,
      readdata => pio_delay_decay_s1_readdata,
      address => pio_delay_decay_s1_address,
      chipselect => pio_delay_decay_s1_chipselect,
      clk => clk_0,
      reset_n => pio_delay_decay_s1_reset_n,
      write_n => pio_delay_decay_s1_write_n,
      writedata => pio_delay_decay_s1_writedata
    );


  --the_pio_delay_length_s1, which is an e_instance
  the_pio_delay_length_s1 : pio_delay_length_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_delay_length_s1 => cpu_data_master_granted_pio_delay_length_s1,
      cpu_data_master_qualified_request_pio_delay_length_s1 => cpu_data_master_qualified_request_pio_delay_length_s1,
      cpu_data_master_read_data_valid_pio_delay_length_s1 => cpu_data_master_read_data_valid_pio_delay_length_s1,
      cpu_data_master_requests_pio_delay_length_s1 => cpu_data_master_requests_pio_delay_length_s1,
      d1_pio_delay_length_s1_end_xfer => d1_pio_delay_length_s1_end_xfer,
      pio_delay_length_s1_address => pio_delay_length_s1_address,
      pio_delay_length_s1_chipselect => pio_delay_length_s1_chipselect,
      pio_delay_length_s1_readdata_from_sa => pio_delay_length_s1_readdata_from_sa,
      pio_delay_length_s1_reset_n => pio_delay_length_s1_reset_n,
      pio_delay_length_s1_write_n => pio_delay_length_s1_write_n,
      pio_delay_length_s1_writedata => pio_delay_length_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_delay_length_s1_readdata => pio_delay_length_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_delay_length, which is an e_ptf_instance
  the_pio_delay_length : pio_delay_length
    port map(
      out_port => internal_out_port_from_the_pio_delay_length,
      readdata => pio_delay_length_s1_readdata,
      address => pio_delay_length_s1_address,
      chipselect => pio_delay_length_s1_chipselect,
      clk => clk_0,
      reset_n => pio_delay_length_s1_reset_n,
      write_n => pio_delay_length_s1_write_n,
      writedata => pio_delay_length_s1_writedata
    );


  --the_pio_master_volume_s1, which is an e_instance
  the_pio_master_volume_s1 : pio_master_volume_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_master_volume_s1 => cpu_data_master_granted_pio_master_volume_s1,
      cpu_data_master_qualified_request_pio_master_volume_s1 => cpu_data_master_qualified_request_pio_master_volume_s1,
      cpu_data_master_read_data_valid_pio_master_volume_s1 => cpu_data_master_read_data_valid_pio_master_volume_s1,
      cpu_data_master_requests_pio_master_volume_s1 => cpu_data_master_requests_pio_master_volume_s1,
      d1_pio_master_volume_s1_end_xfer => d1_pio_master_volume_s1_end_xfer,
      pio_master_volume_s1_address => pio_master_volume_s1_address,
      pio_master_volume_s1_chipselect => pio_master_volume_s1_chipselect,
      pio_master_volume_s1_readdata_from_sa => pio_master_volume_s1_readdata_from_sa,
      pio_master_volume_s1_reset_n => pio_master_volume_s1_reset_n,
      pio_master_volume_s1_write_n => pio_master_volume_s1_write_n,
      pio_master_volume_s1_writedata => pio_master_volume_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_master_volume_s1_readdata => pio_master_volume_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_master_volume, which is an e_ptf_instance
  the_pio_master_volume : pio_master_volume
    port map(
      out_port => internal_out_port_from_the_pio_master_volume,
      readdata => pio_master_volume_s1_readdata,
      address => pio_master_volume_s1_address,
      chipselect => pio_master_volume_s1_chipselect,
      clk => clk_0,
      reset_n => pio_master_volume_s1_reset_n,
      write_n => pio_master_volume_s1_write_n,
      writedata => pio_master_volume_s1_writedata
    );


  --the_pio_octaver_bypass_s1, which is an e_instance
  the_pio_octaver_bypass_s1 : pio_octaver_bypass_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_octaver_bypass_s1 => cpu_data_master_granted_pio_octaver_bypass_s1,
      cpu_data_master_qualified_request_pio_octaver_bypass_s1 => cpu_data_master_qualified_request_pio_octaver_bypass_s1,
      cpu_data_master_read_data_valid_pio_octaver_bypass_s1 => cpu_data_master_read_data_valid_pio_octaver_bypass_s1,
      cpu_data_master_requests_pio_octaver_bypass_s1 => cpu_data_master_requests_pio_octaver_bypass_s1,
      d1_pio_octaver_bypass_s1_end_xfer => d1_pio_octaver_bypass_s1_end_xfer,
      pio_octaver_bypass_s1_address => pio_octaver_bypass_s1_address,
      pio_octaver_bypass_s1_chipselect => pio_octaver_bypass_s1_chipselect,
      pio_octaver_bypass_s1_readdata_from_sa => pio_octaver_bypass_s1_readdata_from_sa,
      pio_octaver_bypass_s1_reset_n => pio_octaver_bypass_s1_reset_n,
      pio_octaver_bypass_s1_write_n => pio_octaver_bypass_s1_write_n,
      pio_octaver_bypass_s1_writedata => pio_octaver_bypass_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_octaver_bypass_s1_readdata => pio_octaver_bypass_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_octaver_bypass, which is an e_ptf_instance
  the_pio_octaver_bypass : pio_octaver_bypass
    port map(
      out_port => internal_out_port_from_the_pio_octaver_bypass,
      readdata => pio_octaver_bypass_s1_readdata,
      address => pio_octaver_bypass_s1_address,
      chipselect => pio_octaver_bypass_s1_chipselect,
      clk => clk_0,
      reset_n => pio_octaver_bypass_s1_reset_n,
      write_n => pio_octaver_bypass_s1_write_n,
      writedata => pio_octaver_bypass_s1_writedata
    );


  --the_pio_octaver_dry_wet_s1, which is an e_instance
  the_pio_octaver_dry_wet_s1 : pio_octaver_dry_wet_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_octaver_dry_wet_s1 => cpu_data_master_granted_pio_octaver_dry_wet_s1,
      cpu_data_master_qualified_request_pio_octaver_dry_wet_s1 => cpu_data_master_qualified_request_pio_octaver_dry_wet_s1,
      cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1 => cpu_data_master_read_data_valid_pio_octaver_dry_wet_s1,
      cpu_data_master_requests_pio_octaver_dry_wet_s1 => cpu_data_master_requests_pio_octaver_dry_wet_s1,
      d1_pio_octaver_dry_wet_s1_end_xfer => d1_pio_octaver_dry_wet_s1_end_xfer,
      pio_octaver_dry_wet_s1_address => pio_octaver_dry_wet_s1_address,
      pio_octaver_dry_wet_s1_chipselect => pio_octaver_dry_wet_s1_chipselect,
      pio_octaver_dry_wet_s1_readdata_from_sa => pio_octaver_dry_wet_s1_readdata_from_sa,
      pio_octaver_dry_wet_s1_reset_n => pio_octaver_dry_wet_s1_reset_n,
      pio_octaver_dry_wet_s1_write_n => pio_octaver_dry_wet_s1_write_n,
      pio_octaver_dry_wet_s1_writedata => pio_octaver_dry_wet_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_octaver_dry_wet_s1_readdata => pio_octaver_dry_wet_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_octaver_dry_wet, which is an e_ptf_instance
  the_pio_octaver_dry_wet : pio_octaver_dry_wet
    port map(
      out_port => internal_out_port_from_the_pio_octaver_dry_wet,
      readdata => pio_octaver_dry_wet_s1_readdata,
      address => pio_octaver_dry_wet_s1_address,
      chipselect => pio_octaver_dry_wet_s1_chipselect,
      clk => clk_0,
      reset_n => pio_octaver_dry_wet_s1_reset_n,
      write_n => pio_octaver_dry_wet_s1_write_n,
      writedata => pio_octaver_dry_wet_s1_writedata
    );


  --the_pio_output_power_left_s1, which is an e_instance
  the_pio_output_power_left_s1 : pio_output_power_left_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_output_power_left_s1 => cpu_data_master_granted_pio_output_power_left_s1,
      cpu_data_master_qualified_request_pio_output_power_left_s1 => cpu_data_master_qualified_request_pio_output_power_left_s1,
      cpu_data_master_read_data_valid_pio_output_power_left_s1 => cpu_data_master_read_data_valid_pio_output_power_left_s1,
      cpu_data_master_requests_pio_output_power_left_s1 => cpu_data_master_requests_pio_output_power_left_s1,
      d1_pio_output_power_left_s1_end_xfer => d1_pio_output_power_left_s1_end_xfer,
      pio_output_power_left_s1_address => pio_output_power_left_s1_address,
      pio_output_power_left_s1_readdata_from_sa => pio_output_power_left_s1_readdata_from_sa,
      pio_output_power_left_s1_reset_n => pio_output_power_left_s1_reset_n,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_write => cpu_data_master_write,
      pio_output_power_left_s1_readdata => pio_output_power_left_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_output_power_left, which is an e_ptf_instance
  the_pio_output_power_left : pio_output_power_left
    port map(
      readdata => pio_output_power_left_s1_readdata,
      address => pio_output_power_left_s1_address,
      clk => clk_0,
      in_port => in_port_to_the_pio_output_power_left,
      reset_n => pio_output_power_left_s1_reset_n
    );


  --the_pio_output_power_right_s1, which is an e_instance
  the_pio_output_power_right_s1 : pio_output_power_right_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_output_power_right_s1 => cpu_data_master_granted_pio_output_power_right_s1,
      cpu_data_master_qualified_request_pio_output_power_right_s1 => cpu_data_master_qualified_request_pio_output_power_right_s1,
      cpu_data_master_read_data_valid_pio_output_power_right_s1 => cpu_data_master_read_data_valid_pio_output_power_right_s1,
      cpu_data_master_requests_pio_output_power_right_s1 => cpu_data_master_requests_pio_output_power_right_s1,
      d1_pio_output_power_right_s1_end_xfer => d1_pio_output_power_right_s1_end_xfer,
      pio_output_power_right_s1_address => pio_output_power_right_s1_address,
      pio_output_power_right_s1_readdata_from_sa => pio_output_power_right_s1_readdata_from_sa,
      pio_output_power_right_s1_reset_n => pio_output_power_right_s1_reset_n,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_write => cpu_data_master_write,
      pio_output_power_right_s1_readdata => pio_output_power_right_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_output_power_right, which is an e_ptf_instance
  the_pio_output_power_right : pio_output_power_right
    port map(
      readdata => pio_output_power_right_s1_readdata,
      address => pio_output_power_right_s1_address,
      clk => clk_0,
      in_port => in_port_to_the_pio_output_power_right,
      reset_n => pio_output_power_right_s1_reset_n
    );


  --the_pio_overdrive_asymmetric_s1, which is an e_instance
  the_pio_overdrive_asymmetric_s1 : pio_overdrive_asymmetric_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_overdrive_asymmetric_s1 => cpu_data_master_granted_pio_overdrive_asymmetric_s1,
      cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1 => cpu_data_master_qualified_request_pio_overdrive_asymmetric_s1,
      cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1 => cpu_data_master_read_data_valid_pio_overdrive_asymmetric_s1,
      cpu_data_master_requests_pio_overdrive_asymmetric_s1 => cpu_data_master_requests_pio_overdrive_asymmetric_s1,
      d1_pio_overdrive_asymmetric_s1_end_xfer => d1_pio_overdrive_asymmetric_s1_end_xfer,
      pio_overdrive_asymmetric_s1_address => pio_overdrive_asymmetric_s1_address,
      pio_overdrive_asymmetric_s1_chipselect => pio_overdrive_asymmetric_s1_chipselect,
      pio_overdrive_asymmetric_s1_readdata_from_sa => pio_overdrive_asymmetric_s1_readdata_from_sa,
      pio_overdrive_asymmetric_s1_reset_n => pio_overdrive_asymmetric_s1_reset_n,
      pio_overdrive_asymmetric_s1_write_n => pio_overdrive_asymmetric_s1_write_n,
      pio_overdrive_asymmetric_s1_writedata => pio_overdrive_asymmetric_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_overdrive_asymmetric_s1_readdata => pio_overdrive_asymmetric_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_overdrive_asymmetric, which is an e_ptf_instance
  the_pio_overdrive_asymmetric : pio_overdrive_asymmetric
    port map(
      out_port => internal_out_port_from_the_pio_overdrive_asymmetric,
      readdata => pio_overdrive_asymmetric_s1_readdata,
      address => pio_overdrive_asymmetric_s1_address,
      chipselect => pio_overdrive_asymmetric_s1_chipselect,
      clk => clk_0,
      reset_n => pio_overdrive_asymmetric_s1_reset_n,
      write_n => pio_overdrive_asymmetric_s1_write_n,
      writedata => pio_overdrive_asymmetric_s1_writedata
    );


  --the_pio_overdrive_bypass_s1, which is an e_instance
  the_pio_overdrive_bypass_s1 : pio_overdrive_bypass_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_overdrive_bypass_s1 => cpu_data_master_granted_pio_overdrive_bypass_s1,
      cpu_data_master_qualified_request_pio_overdrive_bypass_s1 => cpu_data_master_qualified_request_pio_overdrive_bypass_s1,
      cpu_data_master_read_data_valid_pio_overdrive_bypass_s1 => cpu_data_master_read_data_valid_pio_overdrive_bypass_s1,
      cpu_data_master_requests_pio_overdrive_bypass_s1 => cpu_data_master_requests_pio_overdrive_bypass_s1,
      d1_pio_overdrive_bypass_s1_end_xfer => d1_pio_overdrive_bypass_s1_end_xfer,
      pio_overdrive_bypass_s1_address => pio_overdrive_bypass_s1_address,
      pio_overdrive_bypass_s1_chipselect => pio_overdrive_bypass_s1_chipselect,
      pio_overdrive_bypass_s1_readdata_from_sa => pio_overdrive_bypass_s1_readdata_from_sa,
      pio_overdrive_bypass_s1_reset_n => pio_overdrive_bypass_s1_reset_n,
      pio_overdrive_bypass_s1_write_n => pio_overdrive_bypass_s1_write_n,
      pio_overdrive_bypass_s1_writedata => pio_overdrive_bypass_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_overdrive_bypass_s1_readdata => pio_overdrive_bypass_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_overdrive_bypass, which is an e_ptf_instance
  the_pio_overdrive_bypass : pio_overdrive_bypass
    port map(
      out_port => internal_out_port_from_the_pio_overdrive_bypass,
      readdata => pio_overdrive_bypass_s1_readdata,
      address => pio_overdrive_bypass_s1_address,
      chipselect => pio_overdrive_bypass_s1_chipselect,
      clk => clk_0,
      reset_n => pio_overdrive_bypass_s1_reset_n,
      write_n => pio_overdrive_bypass_s1_write_n,
      writedata => pio_overdrive_bypass_s1_writedata
    );


  --the_pio_overdrive_gain_s1, which is an e_instance
  the_pio_overdrive_gain_s1 : pio_overdrive_gain_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_overdrive_gain_s1 => cpu_data_master_granted_pio_overdrive_gain_s1,
      cpu_data_master_qualified_request_pio_overdrive_gain_s1 => cpu_data_master_qualified_request_pio_overdrive_gain_s1,
      cpu_data_master_read_data_valid_pio_overdrive_gain_s1 => cpu_data_master_read_data_valid_pio_overdrive_gain_s1,
      cpu_data_master_requests_pio_overdrive_gain_s1 => cpu_data_master_requests_pio_overdrive_gain_s1,
      d1_pio_overdrive_gain_s1_end_xfer => d1_pio_overdrive_gain_s1_end_xfer,
      pio_overdrive_gain_s1_address => pio_overdrive_gain_s1_address,
      pio_overdrive_gain_s1_chipselect => pio_overdrive_gain_s1_chipselect,
      pio_overdrive_gain_s1_readdata_from_sa => pio_overdrive_gain_s1_readdata_from_sa,
      pio_overdrive_gain_s1_reset_n => pio_overdrive_gain_s1_reset_n,
      pio_overdrive_gain_s1_write_n => pio_overdrive_gain_s1_write_n,
      pio_overdrive_gain_s1_writedata => pio_overdrive_gain_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_overdrive_gain_s1_readdata => pio_overdrive_gain_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_overdrive_gain, which is an e_ptf_instance
  the_pio_overdrive_gain : pio_overdrive_gain
    port map(
      out_port => internal_out_port_from_the_pio_overdrive_gain,
      readdata => pio_overdrive_gain_s1_readdata,
      address => pio_overdrive_gain_s1_address,
      chipselect => pio_overdrive_gain_s1_chipselect,
      clk => clk_0,
      reset_n => pio_overdrive_gain_s1_reset_n,
      write_n => pio_overdrive_gain_s1_write_n,
      writedata => pio_overdrive_gain_s1_writedata
    );


  --the_pio_overdrive_tone_s1, which is an e_instance
  the_pio_overdrive_tone_s1 : pio_overdrive_tone_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_overdrive_tone_s1 => cpu_data_master_granted_pio_overdrive_tone_s1,
      cpu_data_master_qualified_request_pio_overdrive_tone_s1 => cpu_data_master_qualified_request_pio_overdrive_tone_s1,
      cpu_data_master_read_data_valid_pio_overdrive_tone_s1 => cpu_data_master_read_data_valid_pio_overdrive_tone_s1,
      cpu_data_master_requests_pio_overdrive_tone_s1 => cpu_data_master_requests_pio_overdrive_tone_s1,
      d1_pio_overdrive_tone_s1_end_xfer => d1_pio_overdrive_tone_s1_end_xfer,
      pio_overdrive_tone_s1_address => pio_overdrive_tone_s1_address,
      pio_overdrive_tone_s1_chipselect => pio_overdrive_tone_s1_chipselect,
      pio_overdrive_tone_s1_readdata_from_sa => pio_overdrive_tone_s1_readdata_from_sa,
      pio_overdrive_tone_s1_reset_n => pio_overdrive_tone_s1_reset_n,
      pio_overdrive_tone_s1_write_n => pio_overdrive_tone_s1_write_n,
      pio_overdrive_tone_s1_writedata => pio_overdrive_tone_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_overdrive_tone_s1_readdata => pio_overdrive_tone_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_overdrive_tone, which is an e_ptf_instance
  the_pio_overdrive_tone : pio_overdrive_tone
    port map(
      out_port => internal_out_port_from_the_pio_overdrive_tone,
      readdata => pio_overdrive_tone_s1_readdata,
      address => pio_overdrive_tone_s1_address,
      chipselect => pio_overdrive_tone_s1_chipselect,
      clk => clk_0,
      reset_n => pio_overdrive_tone_s1_reset_n,
      write_n => pio_overdrive_tone_s1_write_n,
      writedata => pio_overdrive_tone_s1_writedata
    );


  --the_pio_overdrive_volume_s1, which is an e_instance
  the_pio_overdrive_volume_s1 : pio_overdrive_volume_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_overdrive_volume_s1 => cpu_data_master_granted_pio_overdrive_volume_s1,
      cpu_data_master_qualified_request_pio_overdrive_volume_s1 => cpu_data_master_qualified_request_pio_overdrive_volume_s1,
      cpu_data_master_read_data_valid_pio_overdrive_volume_s1 => cpu_data_master_read_data_valid_pio_overdrive_volume_s1,
      cpu_data_master_requests_pio_overdrive_volume_s1 => cpu_data_master_requests_pio_overdrive_volume_s1,
      d1_pio_overdrive_volume_s1_end_xfer => d1_pio_overdrive_volume_s1_end_xfer,
      pio_overdrive_volume_s1_address => pio_overdrive_volume_s1_address,
      pio_overdrive_volume_s1_chipselect => pio_overdrive_volume_s1_chipselect,
      pio_overdrive_volume_s1_readdata_from_sa => pio_overdrive_volume_s1_readdata_from_sa,
      pio_overdrive_volume_s1_reset_n => pio_overdrive_volume_s1_reset_n,
      pio_overdrive_volume_s1_write_n => pio_overdrive_volume_s1_write_n,
      pio_overdrive_volume_s1_writedata => pio_overdrive_volume_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_overdrive_volume_s1_readdata => pio_overdrive_volume_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_overdrive_volume, which is an e_ptf_instance
  the_pio_overdrive_volume : pio_overdrive_volume
    port map(
      out_port => internal_out_port_from_the_pio_overdrive_volume,
      readdata => pio_overdrive_volume_s1_readdata,
      address => pio_overdrive_volume_s1_address,
      chipselect => pio_overdrive_volume_s1_chipselect,
      clk => clk_0,
      reset_n => pio_overdrive_volume_s1_reset_n,
      write_n => pio_overdrive_volume_s1_write_n,
      writedata => pio_overdrive_volume_s1_writedata
    );


  --the_pio_tremolo_stereo_bypass_s1, which is an e_instance
  the_pio_tremolo_stereo_bypass_s1 : pio_tremolo_stereo_bypass_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_tremolo_stereo_bypass_s1 => cpu_data_master_granted_pio_tremolo_stereo_bypass_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_bypass_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_bypass_s1,
      cpu_data_master_requests_pio_tremolo_stereo_bypass_s1 => cpu_data_master_requests_pio_tremolo_stereo_bypass_s1,
      d1_pio_tremolo_stereo_bypass_s1_end_xfer => d1_pio_tremolo_stereo_bypass_s1_end_xfer,
      pio_tremolo_stereo_bypass_s1_address => pio_tremolo_stereo_bypass_s1_address,
      pio_tremolo_stereo_bypass_s1_chipselect => pio_tremolo_stereo_bypass_s1_chipselect,
      pio_tremolo_stereo_bypass_s1_readdata_from_sa => pio_tremolo_stereo_bypass_s1_readdata_from_sa,
      pio_tremolo_stereo_bypass_s1_reset_n => pio_tremolo_stereo_bypass_s1_reset_n,
      pio_tremolo_stereo_bypass_s1_write_n => pio_tremolo_stereo_bypass_s1_write_n,
      pio_tremolo_stereo_bypass_s1_writedata => pio_tremolo_stereo_bypass_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_tremolo_stereo_bypass_s1_readdata => pio_tremolo_stereo_bypass_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_tremolo_stereo_bypass, which is an e_ptf_instance
  the_pio_tremolo_stereo_bypass : pio_tremolo_stereo_bypass
    port map(
      out_port => internal_out_port_from_the_pio_tremolo_stereo_bypass,
      readdata => pio_tremolo_stereo_bypass_s1_readdata,
      address => pio_tremolo_stereo_bypass_s1_address,
      chipselect => pio_tremolo_stereo_bypass_s1_chipselect,
      clk => clk_0,
      reset_n => pio_tremolo_stereo_bypass_s1_reset_n,
      write_n => pio_tremolo_stereo_bypass_s1_write_n,
      writedata => pio_tremolo_stereo_bypass_s1_writedata
    );


  --the_pio_tremolo_stereo_depth_s1, which is an e_instance
  the_pio_tremolo_stereo_depth_s1 : pio_tremolo_stereo_depth_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_tremolo_stereo_depth_s1 => cpu_data_master_granted_pio_tremolo_stereo_depth_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_depth_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_depth_s1,
      cpu_data_master_requests_pio_tremolo_stereo_depth_s1 => cpu_data_master_requests_pio_tremolo_stereo_depth_s1,
      d1_pio_tremolo_stereo_depth_s1_end_xfer => d1_pio_tremolo_stereo_depth_s1_end_xfer,
      pio_tremolo_stereo_depth_s1_address => pio_tremolo_stereo_depth_s1_address,
      pio_tremolo_stereo_depth_s1_chipselect => pio_tremolo_stereo_depth_s1_chipselect,
      pio_tremolo_stereo_depth_s1_readdata_from_sa => pio_tremolo_stereo_depth_s1_readdata_from_sa,
      pio_tremolo_stereo_depth_s1_reset_n => pio_tremolo_stereo_depth_s1_reset_n,
      pio_tremolo_stereo_depth_s1_write_n => pio_tremolo_stereo_depth_s1_write_n,
      pio_tremolo_stereo_depth_s1_writedata => pio_tremolo_stereo_depth_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_tremolo_stereo_depth_s1_readdata => pio_tremolo_stereo_depth_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_tremolo_stereo_depth, which is an e_ptf_instance
  the_pio_tremolo_stereo_depth : pio_tremolo_stereo_depth
    port map(
      out_port => internal_out_port_from_the_pio_tremolo_stereo_depth,
      readdata => pio_tremolo_stereo_depth_s1_readdata,
      address => pio_tremolo_stereo_depth_s1_address,
      chipselect => pio_tremolo_stereo_depth_s1_chipselect,
      clk => clk_0,
      reset_n => pio_tremolo_stereo_depth_s1_reset_n,
      write_n => pio_tremolo_stereo_depth_s1_write_n,
      writedata => pio_tremolo_stereo_depth_s1_writedata
    );


  --the_pio_tremolo_stereo_mode_s1, which is an e_instance
  the_pio_tremolo_stereo_mode_s1 : pio_tremolo_stereo_mode_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_tremolo_stereo_mode_s1 => cpu_data_master_granted_pio_tremolo_stereo_mode_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_mode_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_mode_s1,
      cpu_data_master_requests_pio_tremolo_stereo_mode_s1 => cpu_data_master_requests_pio_tremolo_stereo_mode_s1,
      d1_pio_tremolo_stereo_mode_s1_end_xfer => d1_pio_tremolo_stereo_mode_s1_end_xfer,
      pio_tremolo_stereo_mode_s1_address => pio_tremolo_stereo_mode_s1_address,
      pio_tremolo_stereo_mode_s1_chipselect => pio_tremolo_stereo_mode_s1_chipselect,
      pio_tremolo_stereo_mode_s1_readdata_from_sa => pio_tremolo_stereo_mode_s1_readdata_from_sa,
      pio_tremolo_stereo_mode_s1_reset_n => pio_tremolo_stereo_mode_s1_reset_n,
      pio_tremolo_stereo_mode_s1_write_n => pio_tremolo_stereo_mode_s1_write_n,
      pio_tremolo_stereo_mode_s1_writedata => pio_tremolo_stereo_mode_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_tremolo_stereo_mode_s1_readdata => pio_tremolo_stereo_mode_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_tremolo_stereo_mode, which is an e_ptf_instance
  the_pio_tremolo_stereo_mode : pio_tremolo_stereo_mode
    port map(
      out_port => internal_out_port_from_the_pio_tremolo_stereo_mode,
      readdata => pio_tremolo_stereo_mode_s1_readdata,
      address => pio_tremolo_stereo_mode_s1_address,
      chipselect => pio_tremolo_stereo_mode_s1_chipselect,
      clk => clk_0,
      reset_n => pio_tremolo_stereo_mode_s1_reset_n,
      write_n => pio_tremolo_stereo_mode_s1_write_n,
      writedata => pio_tremolo_stereo_mode_s1_writedata
    );


  --the_pio_tremolo_stereo_sweep_a_s1, which is an e_instance
  the_pio_tremolo_stereo_sweep_a_s1 : pio_tremolo_stereo_sweep_a_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_granted_pio_tremolo_stereo_sweep_a_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_a_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_a_s1,
      cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1 => cpu_data_master_requests_pio_tremolo_stereo_sweep_a_s1,
      d1_pio_tremolo_stereo_sweep_a_s1_end_xfer => d1_pio_tremolo_stereo_sweep_a_s1_end_xfer,
      pio_tremolo_stereo_sweep_a_s1_address => pio_tremolo_stereo_sweep_a_s1_address,
      pio_tremolo_stereo_sweep_a_s1_chipselect => pio_tremolo_stereo_sweep_a_s1_chipselect,
      pio_tremolo_stereo_sweep_a_s1_readdata_from_sa => pio_tremolo_stereo_sweep_a_s1_readdata_from_sa,
      pio_tremolo_stereo_sweep_a_s1_reset_n => pio_tremolo_stereo_sweep_a_s1_reset_n,
      pio_tremolo_stereo_sweep_a_s1_write_n => pio_tremolo_stereo_sweep_a_s1_write_n,
      pio_tremolo_stereo_sweep_a_s1_writedata => pio_tremolo_stereo_sweep_a_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_tremolo_stereo_sweep_a_s1_readdata => pio_tremolo_stereo_sweep_a_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_tremolo_stereo_sweep_a, which is an e_ptf_instance
  the_pio_tremolo_stereo_sweep_a : pio_tremolo_stereo_sweep_a
    port map(
      out_port => internal_out_port_from_the_pio_tremolo_stereo_sweep_a,
      readdata => pio_tremolo_stereo_sweep_a_s1_readdata,
      address => pio_tremolo_stereo_sweep_a_s1_address,
      chipselect => pio_tremolo_stereo_sweep_a_s1_chipselect,
      clk => clk_0,
      reset_n => pio_tremolo_stereo_sweep_a_s1_reset_n,
      write_n => pio_tremolo_stereo_sweep_a_s1_write_n,
      writedata => pio_tremolo_stereo_sweep_a_s1_writedata
    );


  --the_pio_tremolo_stereo_sweep_b_s1, which is an e_instance
  the_pio_tremolo_stereo_sweep_b_s1 : pio_tremolo_stereo_sweep_b_s1_arbitrator
    port map(
      cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_granted_pio_tremolo_stereo_sweep_b_s1,
      cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_qualified_request_pio_tremolo_stereo_sweep_b_s1,
      cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_read_data_valid_pio_tremolo_stereo_sweep_b_s1,
      cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1 => cpu_data_master_requests_pio_tremolo_stereo_sweep_b_s1,
      d1_pio_tremolo_stereo_sweep_b_s1_end_xfer => d1_pio_tremolo_stereo_sweep_b_s1_end_xfer,
      pio_tremolo_stereo_sweep_b_s1_address => pio_tremolo_stereo_sweep_b_s1_address,
      pio_tremolo_stereo_sweep_b_s1_chipselect => pio_tremolo_stereo_sweep_b_s1_chipselect,
      pio_tremolo_stereo_sweep_b_s1_readdata_from_sa => pio_tremolo_stereo_sweep_b_s1_readdata_from_sa,
      pio_tremolo_stereo_sweep_b_s1_reset_n => pio_tremolo_stereo_sweep_b_s1_reset_n,
      pio_tremolo_stereo_sweep_b_s1_write_n => pio_tremolo_stereo_sweep_b_s1_write_n,
      pio_tremolo_stereo_sweep_b_s1_writedata => pio_tremolo_stereo_sweep_b_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pio_tremolo_stereo_sweep_b_s1_readdata => pio_tremolo_stereo_sweep_b_s1_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pio_tremolo_stereo_sweep_b, which is an e_ptf_instance
  the_pio_tremolo_stereo_sweep_b : pio_tremolo_stereo_sweep_b
    port map(
      out_port => internal_out_port_from_the_pio_tremolo_stereo_sweep_b,
      readdata => pio_tremolo_stereo_sweep_b_s1_readdata,
      address => pio_tremolo_stereo_sweep_b_s1_address,
      chipselect => pio_tremolo_stereo_sweep_b_s1_chipselect,
      clk => clk_0,
      reset_n => pio_tremolo_stereo_sweep_b_s1_reset_n,
      write_n => pio_tremolo_stereo_sweep_b_s1_write_n,
      writedata => pio_tremolo_stereo_sweep_b_s1_writedata
    );


  --the_pixel_buffer_avalon_pixel_buffer_slave, which is an e_instance
  the_pixel_buffer_avalon_pixel_buffer_slave : pixel_buffer_avalon_pixel_buffer_slave_arbitrator
    port map(
      cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_granted_pixel_buffer_avalon_pixel_buffer_slave,
      cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_qualified_request_pixel_buffer_avalon_pixel_buffer_slave,
      cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave,
      cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave => cpu_data_master_requests_pixel_buffer_avalon_pixel_buffer_slave,
      d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer => d1_pixel_buffer_avalon_pixel_buffer_slave_end_xfer,
      pixel_buffer_avalon_pixel_buffer_slave_address => pixel_buffer_avalon_pixel_buffer_slave_address,
      pixel_buffer_avalon_pixel_buffer_slave_byteenable => pixel_buffer_avalon_pixel_buffer_slave_byteenable,
      pixel_buffer_avalon_pixel_buffer_slave_read => pixel_buffer_avalon_pixel_buffer_slave_read,
      pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa => pixel_buffer_avalon_pixel_buffer_slave_readdata_from_sa,
      pixel_buffer_avalon_pixel_buffer_slave_reset => pixel_buffer_avalon_pixel_buffer_slave_reset,
      pixel_buffer_avalon_pixel_buffer_slave_write => pixel_buffer_avalon_pixel_buffer_slave_write,
      pixel_buffer_avalon_pixel_buffer_slave_writedata => pixel_buffer_avalon_pixel_buffer_slave_writedata,
      registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave => registered_cpu_data_master_read_data_valid_pixel_buffer_avalon_pixel_buffer_slave,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      pixel_buffer_avalon_pixel_buffer_slave_readdata => pixel_buffer_avalon_pixel_buffer_slave_readdata,
      reset_n => clk_0_reset_n
    );


  --the_pixel_buffer_avalon_pixel_buffer_master, which is an e_instance
  the_pixel_buffer_avalon_pixel_buffer_master : pixel_buffer_avalon_pixel_buffer_master_arbitrator
    port map(
      pixel_buffer_avalon_pixel_buffer_master_address_to_slave => pixel_buffer_avalon_pixel_buffer_master_address_to_slave,
      pixel_buffer_avalon_pixel_buffer_master_latency_counter => pixel_buffer_avalon_pixel_buffer_master_latency_counter,
      pixel_buffer_avalon_pixel_buffer_master_readdata => pixel_buffer_avalon_pixel_buffer_master_readdata,
      pixel_buffer_avalon_pixel_buffer_master_readdatavalid => pixel_buffer_avalon_pixel_buffer_master_readdatavalid,
      pixel_buffer_avalon_pixel_buffer_master_waitrequest => pixel_buffer_avalon_pixel_buffer_master_waitrequest,
      clk => clk_0,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      pixel_buffer_avalon_pixel_buffer_master_address => pixel_buffer_avalon_pixel_buffer_master_address,
      pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1,
      pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1,
      pixel_buffer_avalon_pixel_buffer_master_read => pixel_buffer_avalon_pixel_buffer_master_read,
      pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1,
      pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register => pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register,
      pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1,
      reset_n => clk_0_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa
    );


  --the_pixel_buffer_avalon_pixel_buffer_source, which is an e_instance
  the_pixel_buffer_avalon_pixel_buffer_source : pixel_buffer_avalon_pixel_buffer_source_arbitrator
    port map(
      pixel_buffer_avalon_pixel_buffer_source_ready => pixel_buffer_avalon_pixel_buffer_source_ready,
      alpha_blending_avalon_background_sink_ready_from_sa => alpha_blending_avalon_background_sink_ready_from_sa,
      clk => clk_0,
      pixel_buffer_avalon_pixel_buffer_source_data => pixel_buffer_avalon_pixel_buffer_source_data,
      pixel_buffer_avalon_pixel_buffer_source_empty => pixel_buffer_avalon_pixel_buffer_source_empty,
      pixel_buffer_avalon_pixel_buffer_source_endofpacket => pixel_buffer_avalon_pixel_buffer_source_endofpacket,
      pixel_buffer_avalon_pixel_buffer_source_startofpacket => pixel_buffer_avalon_pixel_buffer_source_startofpacket,
      pixel_buffer_avalon_pixel_buffer_source_valid => pixel_buffer_avalon_pixel_buffer_source_valid,
      reset_n => clk_0_reset_n
    );


  --the_pixel_buffer, which is an e_ptf_instance
  the_pixel_buffer : pixel_buffer
    port map(
      master_address => pixel_buffer_avalon_pixel_buffer_master_address,
      master_arbiterlock => pixel_buffer_avalon_pixel_buffer_master_arbiterlock,
      master_read => pixel_buffer_avalon_pixel_buffer_master_read,
      slave_readdata => pixel_buffer_avalon_pixel_buffer_slave_readdata,
      stream_data => pixel_buffer_avalon_pixel_buffer_source_data,
      stream_empty => pixel_buffer_avalon_pixel_buffer_source_empty,
      stream_endofpacket => pixel_buffer_avalon_pixel_buffer_source_endofpacket,
      stream_startofpacket => pixel_buffer_avalon_pixel_buffer_source_startofpacket,
      stream_valid => pixel_buffer_avalon_pixel_buffer_source_valid,
      clk => clk_0,
      master_readdata => pixel_buffer_avalon_pixel_buffer_master_readdata,
      master_readdatavalid => pixel_buffer_avalon_pixel_buffer_master_readdatavalid,
      master_waitrequest => pixel_buffer_avalon_pixel_buffer_master_waitrequest,
      reset => pixel_buffer_avalon_pixel_buffer_slave_reset,
      slave_address => pixel_buffer_avalon_pixel_buffer_slave_address,
      slave_byteenable => pixel_buffer_avalon_pixel_buffer_slave_byteenable,
      slave_read => pixel_buffer_avalon_pixel_buffer_slave_read,
      slave_write => pixel_buffer_avalon_pixel_buffer_slave_write,
      slave_writedata => pixel_buffer_avalon_pixel_buffer_slave_writedata,
      stream_ready => pixel_buffer_avalon_pixel_buffer_source_ready
    );


  --the_ps2_avalon_ps2_slave, which is an e_instance
  the_ps2_avalon_ps2_slave : ps2_avalon_ps2_slave_arbitrator
    port map(
      cpu_data_master_granted_ps2_avalon_ps2_slave => cpu_data_master_granted_ps2_avalon_ps2_slave,
      cpu_data_master_qualified_request_ps2_avalon_ps2_slave => cpu_data_master_qualified_request_ps2_avalon_ps2_slave,
      cpu_data_master_read_data_valid_ps2_avalon_ps2_slave => cpu_data_master_read_data_valid_ps2_avalon_ps2_slave,
      cpu_data_master_requests_ps2_avalon_ps2_slave => cpu_data_master_requests_ps2_avalon_ps2_slave,
      d1_ps2_avalon_ps2_slave_end_xfer => d1_ps2_avalon_ps2_slave_end_xfer,
      ps2_avalon_ps2_slave_address => ps2_avalon_ps2_slave_address,
      ps2_avalon_ps2_slave_byteenable => ps2_avalon_ps2_slave_byteenable,
      ps2_avalon_ps2_slave_chipselect => ps2_avalon_ps2_slave_chipselect,
      ps2_avalon_ps2_slave_irq_from_sa => ps2_avalon_ps2_slave_irq_from_sa,
      ps2_avalon_ps2_slave_read => ps2_avalon_ps2_slave_read,
      ps2_avalon_ps2_slave_readdata_from_sa => ps2_avalon_ps2_slave_readdata_from_sa,
      ps2_avalon_ps2_slave_reset => ps2_avalon_ps2_slave_reset,
      ps2_avalon_ps2_slave_waitrequest_from_sa => ps2_avalon_ps2_slave_waitrequest_from_sa,
      ps2_avalon_ps2_slave_write => ps2_avalon_ps2_slave_write,
      ps2_avalon_ps2_slave_writedata => ps2_avalon_ps2_slave_writedata,
      registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave => registered_cpu_data_master_read_data_valid_ps2_avalon_ps2_slave,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      ps2_avalon_ps2_slave_irq => ps2_avalon_ps2_slave_irq,
      ps2_avalon_ps2_slave_readdata => ps2_avalon_ps2_slave_readdata,
      ps2_avalon_ps2_slave_waitrequest => ps2_avalon_ps2_slave_waitrequest,
      reset_n => clk_0_reset_n
    );


  --the_ps2, which is an e_ptf_instance
  the_ps2 : ps2
    port map(
      PS2_CLK => PS2_CLK_to_and_from_the_ps2,
      PS2_DAT => PS2_DAT_to_and_from_the_ps2,
      irq => ps2_avalon_ps2_slave_irq,
      readdata => ps2_avalon_ps2_slave_readdata,
      waitrequest => ps2_avalon_ps2_slave_waitrequest,
      address => ps2_avalon_ps2_slave_address,
      byteenable => ps2_avalon_ps2_slave_byteenable,
      chipselect => ps2_avalon_ps2_slave_chipselect,
      clk => clk_0,
      read => ps2_avalon_ps2_slave_read,
      reset => ps2_avalon_ps2_slave_reset,
      write => ps2_avalon_ps2_slave_write,
      writedata => ps2_avalon_ps2_slave_writedata
    );


  --the_sdram_s1, which is an e_instance
  the_sdram_s1 : sdram_s1_arbitrator
    port map(
      cpu_data_master_byteenable_sdram_s1 => cpu_data_master_byteenable_sdram_s1,
      cpu_data_master_granted_sdram_s1 => cpu_data_master_granted_sdram_s1,
      cpu_data_master_qualified_request_sdram_s1 => cpu_data_master_qualified_request_sdram_s1,
      cpu_data_master_read_data_valid_sdram_s1 => cpu_data_master_read_data_valid_sdram_s1,
      cpu_data_master_read_data_valid_sdram_s1_shift_register => cpu_data_master_read_data_valid_sdram_s1_shift_register,
      cpu_data_master_requests_sdram_s1 => cpu_data_master_requests_sdram_s1,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      membuffer_0_byteenable_sdram_s1 => membuffer_0_byteenable_sdram_s1,
      membuffer_0_granted_sdram_s1 => membuffer_0_granted_sdram_s1,
      membuffer_0_qualified_request_sdram_s1 => membuffer_0_qualified_request_sdram_s1,
      membuffer_0_read_data_valid_sdram_s1 => membuffer_0_read_data_valid_sdram_s1,
      membuffer_0_read_data_valid_sdram_s1_shift_register => membuffer_0_read_data_valid_sdram_s1_shift_register,
      membuffer_0_requests_sdram_s1 => membuffer_0_requests_sdram_s1,
      pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_granted_sdram_s1,
      pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_qualified_request_sdram_s1,
      pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1,
      pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register => pixel_buffer_avalon_pixel_buffer_master_read_data_valid_sdram_s1_shift_register,
      pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1 => pixel_buffer_avalon_pixel_buffer_master_requests_sdram_s1,
      sdram_s1_address => sdram_s1_address,
      sdram_s1_byteenable_n => sdram_s1_byteenable_n,
      sdram_s1_chipselect => sdram_s1_chipselect,
      sdram_s1_read_n => sdram_s1_read_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_reset_n => sdram_s1_reset_n,
      sdram_s1_waitrequest_from_sa => sdram_s1_waitrequest_from_sa,
      sdram_s1_write_n => sdram_s1_write_n,
      sdram_s1_writedata => sdram_s1_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_16 => cpu_data_master_dbs_write_16,
      cpu_data_master_no_byte_enables_and_last_term => cpu_data_master_no_byte_enables_and_last_term,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      membuffer_0_avalon_master_address_to_slave => membuffer_0_avalon_master_address_to_slave,
      membuffer_0_avalon_master_read => membuffer_0_avalon_master_read,
      membuffer_0_avalon_master_write => membuffer_0_avalon_master_write,
      membuffer_0_dbs_address => membuffer_0_dbs_address,
      membuffer_0_dbs_write_16 => membuffer_0_dbs_write_16,
      pixel_buffer_avalon_pixel_buffer_master_address_to_slave => pixel_buffer_avalon_pixel_buffer_master_address_to_slave,
      pixel_buffer_avalon_pixel_buffer_master_arbiterlock => pixel_buffer_avalon_pixel_buffer_master_arbiterlock,
      pixel_buffer_avalon_pixel_buffer_master_latency_counter => pixel_buffer_avalon_pixel_buffer_master_latency_counter,
      pixel_buffer_avalon_pixel_buffer_master_read => pixel_buffer_avalon_pixel_buffer_master_read,
      reset_n => clk_0_reset_n,
      sdram_s1_readdata => sdram_s1_readdata,
      sdram_s1_readdatavalid => sdram_s1_readdatavalid,
      sdram_s1_waitrequest => sdram_s1_waitrequest
    );


  --the_sdram, which is an e_ptf_instance
  the_sdram : sdram
    port map(
      za_data => sdram_s1_readdata,
      za_valid => sdram_s1_readdatavalid,
      za_waitrequest => sdram_s1_waitrequest,
      zs_addr => internal_zs_addr_from_the_sdram,
      zs_ba => internal_zs_ba_from_the_sdram,
      zs_cas_n => internal_zs_cas_n_from_the_sdram,
      zs_cke => internal_zs_cke_from_the_sdram,
      zs_cs_n => internal_zs_cs_n_from_the_sdram,
      zs_dq => zs_dq_to_and_from_the_sdram,
      zs_dqm => internal_zs_dqm_from_the_sdram,
      zs_ras_n => internal_zs_ras_n_from_the_sdram,
      zs_we_n => internal_zs_we_n_from_the_sdram,
      az_addr => sdram_s1_address,
      az_be_n => sdram_s1_byteenable_n,
      az_cs => sdram_s1_chipselect,
      az_data => sdram_s1_writedata,
      az_rd_n => sdram_s1_read_n,
      az_wr_n => sdram_s1_write_n,
      clk => clk_0,
      reset_n => sdram_s1_reset_n
    );


  --the_sram_avalon_sram_slave, which is an e_instance
  the_sram_avalon_sram_slave : sram_avalon_sram_slave_arbitrator
    port map(
      cpu_data_master_byteenable_sram_avalon_sram_slave => cpu_data_master_byteenable_sram_avalon_sram_slave,
      cpu_data_master_granted_sram_avalon_sram_slave => cpu_data_master_granted_sram_avalon_sram_slave,
      cpu_data_master_qualified_request_sram_avalon_sram_slave => cpu_data_master_qualified_request_sram_avalon_sram_slave,
      cpu_data_master_read_data_valid_sram_avalon_sram_slave => cpu_data_master_read_data_valid_sram_avalon_sram_slave,
      cpu_data_master_requests_sram_avalon_sram_slave => cpu_data_master_requests_sram_avalon_sram_slave,
      cpu_instruction_master_granted_sram_avalon_sram_slave => cpu_instruction_master_granted_sram_avalon_sram_slave,
      cpu_instruction_master_qualified_request_sram_avalon_sram_slave => cpu_instruction_master_qualified_request_sram_avalon_sram_slave,
      cpu_instruction_master_read_data_valid_sram_avalon_sram_slave => cpu_instruction_master_read_data_valid_sram_avalon_sram_slave,
      cpu_instruction_master_requests_sram_avalon_sram_slave => cpu_instruction_master_requests_sram_avalon_sram_slave,
      d1_sram_avalon_sram_slave_end_xfer => d1_sram_avalon_sram_slave_end_xfer,
      registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave => registered_cpu_data_master_read_data_valid_sram_avalon_sram_slave,
      sram_avalon_sram_slave_address => sram_avalon_sram_slave_address,
      sram_avalon_sram_slave_byteenable => sram_avalon_sram_slave_byteenable,
      sram_avalon_sram_slave_read => sram_avalon_sram_slave_read,
      sram_avalon_sram_slave_readdata_from_sa => sram_avalon_sram_slave_readdata_from_sa,
      sram_avalon_sram_slave_reset => sram_avalon_sram_slave_reset,
      sram_avalon_sram_slave_write => sram_avalon_sram_slave_write,
      sram_avalon_sram_slave_writedata => sram_avalon_sram_slave_writedata,
      clk => clk_0,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_dbs_address => cpu_data_master_dbs_address,
      cpu_data_master_dbs_write_16 => cpu_data_master_dbs_write_16,
      cpu_data_master_no_byte_enables_and_last_term => cpu_data_master_no_byte_enables_and_last_term,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      cpu_data_master_write => cpu_data_master_write,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_dbs_address => cpu_instruction_master_dbs_address,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      reset_n => clk_0_reset_n,
      sram_avalon_sram_slave_readdata => sram_avalon_sram_slave_readdata
    );


  --the_sram, which is an e_ptf_instance
  the_sram : sram
    port map(
      SRAM_ADDR => internal_SRAM_ADDR_from_the_sram,
      SRAM_CE_N => internal_SRAM_CE_N_from_the_sram,
      SRAM_DQ => SRAM_DQ_to_and_from_the_sram,
      SRAM_LB_N => internal_SRAM_LB_N_from_the_sram,
      SRAM_OE_N => internal_SRAM_OE_N_from_the_sram,
      SRAM_UB_N => internal_SRAM_UB_N_from_the_sram,
      SRAM_WE_N => internal_SRAM_WE_N_from_the_sram,
      readdata => sram_avalon_sram_slave_readdata,
      address => sram_avalon_sram_slave_address,
      byteenable => sram_avalon_sram_slave_byteenable,
      clk => clk_0,
      read => sram_avalon_sram_slave_read,
      reset => sram_avalon_sram_slave_reset,
      write => sram_avalon_sram_slave_write,
      writedata => sram_avalon_sram_slave_writedata
    );


  --the_vga_avalon_vga_sink, which is an e_instance
  the_vga_avalon_vga_sink : vga_avalon_vga_sink_arbitrator
    port map(
      vga_avalon_vga_sink_data => vga_avalon_vga_sink_data,
      vga_avalon_vga_sink_empty => vga_avalon_vga_sink_empty,
      vga_avalon_vga_sink_endofpacket => vga_avalon_vga_sink_endofpacket,
      vga_avalon_vga_sink_ready_from_sa => vga_avalon_vga_sink_ready_from_sa,
      vga_avalon_vga_sink_reset => vga_avalon_vga_sink_reset,
      vga_avalon_vga_sink_startofpacket => vga_avalon_vga_sink_startofpacket,
      vga_avalon_vga_sink_valid => vga_avalon_vga_sink_valid,
      alpha_blending_avalon_blended_source_data => alpha_blending_avalon_blended_source_data,
      alpha_blending_avalon_blended_source_empty => alpha_blending_avalon_blended_source_empty,
      alpha_blending_avalon_blended_source_endofpacket => alpha_blending_avalon_blended_source_endofpacket,
      alpha_blending_avalon_blended_source_startofpacket => alpha_blending_avalon_blended_source_startofpacket,
      alpha_blending_avalon_blended_source_valid => alpha_blending_avalon_blended_source_valid,
      clk => clk_0,
      reset_n => clk_0_reset_n,
      vga_avalon_vga_sink_ready => vga_avalon_vga_sink_ready
    );


  --the_vga, which is an e_ptf_instance
  the_vga : vga
    port map(
      VGA_B => internal_VGA_B_from_the_vga,
      VGA_BLANK => internal_VGA_BLANK_from_the_vga,
      VGA_G => internal_VGA_G_from_the_vga,
      VGA_HS => internal_VGA_HS_from_the_vga,
      VGA_R => internal_VGA_R_from_the_vga,
      VGA_SYNC => internal_VGA_SYNC_from_the_vga,
      VGA_VS => internal_VGA_VS_from_the_vga,
      ready => vga_avalon_vga_sink_ready,
      clk => clk_0,
      data => vga_avalon_vga_sink_data,
      empty => vga_avalon_vga_sink_empty,
      endofpacket => vga_avalon_vga_sink_endofpacket,
      reset => vga_avalon_vga_sink_reset,
      startofpacket => vga_avalon_vga_sink_startofpacket,
      valid => vga_avalon_vga_sink_valid
    );


  --reset is asserted asynchronously and deasserted synchronously
  VGAProc_reset_clk_0_domain_synch : VGAProc_reset_clk_0_domain_synch_module
    port map(
      data_out => clk_0_reset_n,
      clk => clk_0,
      data_in => module_input9,
      reset_n => reset_n_sources
    );

  module_input9 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_resetrequest_from_sa))))));
  --vhdl renameroo for output signals
  FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 <= internal_FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0;
  --vhdl renameroo for output signals
  FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 <= internal_FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0;
  --vhdl renameroo for output signals
  FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 <= internal_FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0;
  --vhdl renameroo for output signals
  FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 <= internal_FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0;
  --vhdl renameroo for output signals
  FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 <= internal_FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0;
  --vhdl renameroo for output signals
  I2C_SCLK_from_the_audio_and_video_config_0 <= internal_I2C_SCLK_from_the_audio_and_video_config_0;
  --vhdl renameroo for output signals
  SRAM_ADDR_from_the_sram <= internal_SRAM_ADDR_from_the_sram;
  --vhdl renameroo for output signals
  SRAM_CE_N_from_the_sram <= internal_SRAM_CE_N_from_the_sram;
  --vhdl renameroo for output signals
  SRAM_LB_N_from_the_sram <= internal_SRAM_LB_N_from_the_sram;
  --vhdl renameroo for output signals
  SRAM_OE_N_from_the_sram <= internal_SRAM_OE_N_from_the_sram;
  --vhdl renameroo for output signals
  SRAM_UB_N_from_the_sram <= internal_SRAM_UB_N_from_the_sram;
  --vhdl renameroo for output signals
  SRAM_WE_N_from_the_sram <= internal_SRAM_WE_N_from_the_sram;
  --vhdl renameroo for output signals
  VGA_BLANK_from_the_vga <= internal_VGA_BLANK_from_the_vga;
  --vhdl renameroo for output signals
  VGA_B_from_the_vga <= internal_VGA_B_from_the_vga;
  --vhdl renameroo for output signals
  VGA_G_from_the_vga <= internal_VGA_G_from_the_vga;
  --vhdl renameroo for output signals
  VGA_HS_from_the_vga <= internal_VGA_HS_from_the_vga;
  --vhdl renameroo for output signals
  VGA_R_from_the_vga <= internal_VGA_R_from_the_vga;
  --vhdl renameroo for output signals
  VGA_SYNC_from_the_vga <= internal_VGA_SYNC_from_the_vga;
  --vhdl renameroo for output signals
  VGA_VS_from_the_vga <= internal_VGA_VS_from_the_vga;
  --vhdl renameroo for output signals
  out_port_from_the_pio_bitcrusher_bypass <= internal_out_port_from_the_pio_bitcrusher_bypass;
  --vhdl renameroo for output signals
  out_port_from_the_pio_bitcrusher_crush <= internal_out_port_from_the_pio_bitcrusher_crush;
  --vhdl renameroo for output signals
  out_port_from_the_pio_bitcrusher_downsample <= internal_out_port_from_the_pio_bitcrusher_downsample;
  --vhdl renameroo for output signals
  out_port_from_the_pio_bitcrusher_drywet <= internal_out_port_from_the_pio_bitcrusher_drywet;
  --vhdl renameroo for output signals
  out_port_from_the_pio_bitcrusher_flavor <= internal_out_port_from_the_pio_bitcrusher_flavor;
  --vhdl renameroo for output signals
  out_port_from_the_pio_bitcrusher_tone <= internal_out_port_from_the_pio_bitcrusher_tone;
  --vhdl renameroo for output signals
  out_port_from_the_pio_compressor_bypass <= internal_out_port_from_the_pio_compressor_bypass;
  --vhdl renameroo for output signals
  out_port_from_the_pio_compressor_gain <= internal_out_port_from_the_pio_compressor_gain;
  --vhdl renameroo for output signals
  out_port_from_the_pio_compressor_treshold <= internal_out_port_from_the_pio_compressor_treshold;
  --vhdl renameroo for output signals
  out_port_from_the_pio_delay_bypass <= internal_out_port_from_the_pio_delay_bypass;
  --vhdl renameroo for output signals
  out_port_from_the_pio_delay_decay <= internal_out_port_from_the_pio_delay_decay;
  --vhdl renameroo for output signals
  out_port_from_the_pio_delay_length <= internal_out_port_from_the_pio_delay_length;
  --vhdl renameroo for output signals
  out_port_from_the_pio_master_volume <= internal_out_port_from_the_pio_master_volume;
  --vhdl renameroo for output signals
  out_port_from_the_pio_octaver_bypass <= internal_out_port_from_the_pio_octaver_bypass;
  --vhdl renameroo for output signals
  out_port_from_the_pio_octaver_dry_wet <= internal_out_port_from_the_pio_octaver_dry_wet;
  --vhdl renameroo for output signals
  out_port_from_the_pio_overdrive_asymmetric <= internal_out_port_from_the_pio_overdrive_asymmetric;
  --vhdl renameroo for output signals
  out_port_from_the_pio_overdrive_bypass <= internal_out_port_from_the_pio_overdrive_bypass;
  --vhdl renameroo for output signals
  out_port_from_the_pio_overdrive_gain <= internal_out_port_from_the_pio_overdrive_gain;
  --vhdl renameroo for output signals
  out_port_from_the_pio_overdrive_tone <= internal_out_port_from_the_pio_overdrive_tone;
  --vhdl renameroo for output signals
  out_port_from_the_pio_overdrive_volume <= internal_out_port_from_the_pio_overdrive_volume;
  --vhdl renameroo for output signals
  out_port_from_the_pio_tremolo_stereo_bypass <= internal_out_port_from_the_pio_tremolo_stereo_bypass;
  --vhdl renameroo for output signals
  out_port_from_the_pio_tremolo_stereo_depth <= internal_out_port_from_the_pio_tremolo_stereo_depth;
  --vhdl renameroo for output signals
  out_port_from_the_pio_tremolo_stereo_mode <= internal_out_port_from_the_pio_tremolo_stereo_mode;
  --vhdl renameroo for output signals
  out_port_from_the_pio_tremolo_stereo_sweep_a <= internal_out_port_from_the_pio_tremolo_stereo_sweep_a;
  --vhdl renameroo for output signals
  out_port_from_the_pio_tremolo_stereo_sweep_b <= internal_out_port_from_the_pio_tremolo_stereo_sweep_b;
  --vhdl renameroo for output signals
  sample_left_out_from_the_membuffer_0 <= internal_sample_left_out_from_the_membuffer_0;
  --vhdl renameroo for output signals
  sample_right_out_from_the_membuffer_0 <= internal_sample_right_out_from_the_membuffer_0;
  --vhdl renameroo for output signals
  zs_addr_from_the_sdram <= internal_zs_addr_from_the_sdram;
  --vhdl renameroo for output signals
  zs_ba_from_the_sdram <= internal_zs_ba_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cas_n_from_the_sdram <= internal_zs_cas_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cke_from_the_sdram <= internal_zs_cke_from_the_sdram;
  --vhdl renameroo for output signals
  zs_cs_n_from_the_sdram <= internal_zs_cs_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_dqm_from_the_sdram <= internal_zs_dqm_from_the_sdram;
  --vhdl renameroo for output signals
  zs_ras_n_from_the_sdram <= internal_zs_ras_n_from_the_sdram;
  --vhdl renameroo for output signals
  zs_we_n_from_the_sdram <= internal_zs_we_n_from_the_sdram;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component VGAProc is 
           port (
                 -- 1) global signals:
                    signal clk_0 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0
                    signal FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;
                    signal FL_DQ_to_and_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;
                    signal FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;
                    signal FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 : OUT STD_LOGIC;

                 -- the_analyzer_input_left
                    signal x_in_to_the_analyzer_input_left : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal y_in_to_the_analyzer_input_left : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

                 -- the_analyzer_input_right
                    signal x_in_to_the_analyzer_input_right : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal y_in_to_the_analyzer_input_right : IN STD_LOGIC_VECTOR (63 DOWNTO 0);

                 -- the_audio_and_video_config_0
                    signal I2C_SCLK_from_the_audio_and_video_config_0 : OUT STD_LOGIC;
                    signal I2C_SDAT_to_and_from_the_audio_and_video_config_0 : INOUT STD_LOGIC;

                 -- the_membuffer_0
                    signal delay_time_to_the_membuffer_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sample_clk_to_the_membuffer_0 : IN STD_LOGIC;
                    signal sample_left_in_to_the_membuffer_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sample_left_out_from_the_membuffer_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sample_right_in_to_the_membuffer_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sample_right_out_from_the_membuffer_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_bitcrusher_bypass
                    signal out_port_from_the_pio_bitcrusher_bypass : OUT STD_LOGIC;

                 -- the_pio_bitcrusher_crush
                    signal out_port_from_the_pio_bitcrusher_crush : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_pio_bitcrusher_downsample
                    signal out_port_from_the_pio_bitcrusher_downsample : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_pio_bitcrusher_drywet
                    signal out_port_from_the_pio_bitcrusher_drywet : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_bitcrusher_flavor
                    signal out_port_from_the_pio_bitcrusher_flavor : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_pio_bitcrusher_tone
                    signal out_port_from_the_pio_bitcrusher_tone : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_compressor_bypass
                    signal out_port_from_the_pio_compressor_bypass : OUT STD_LOGIC;

                 -- the_pio_compressor_gain
                    signal out_port_from_the_pio_compressor_gain : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_pio_compressor_treshold
                    signal out_port_from_the_pio_compressor_treshold : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_delay_bypass
                    signal out_port_from_the_pio_delay_bypass : OUT STD_LOGIC;

                 -- the_pio_delay_decay
                    signal out_port_from_the_pio_delay_decay : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_pio_delay_length
                    signal out_port_from_the_pio_delay_length : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_master_volume
                    signal out_port_from_the_pio_master_volume : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_octaver_bypass
                    signal out_port_from_the_pio_octaver_bypass : OUT STD_LOGIC;

                 -- the_pio_octaver_dry_wet
                    signal out_port_from_the_pio_octaver_dry_wet : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_output_power_left
                    signal in_port_to_the_pio_output_power_left : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_output_power_right
                    signal in_port_to_the_pio_output_power_right : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_overdrive_asymmetric
                    signal out_port_from_the_pio_overdrive_asymmetric : OUT STD_LOGIC;

                 -- the_pio_overdrive_bypass
                    signal out_port_from_the_pio_overdrive_bypass : OUT STD_LOGIC;

                 -- the_pio_overdrive_gain
                    signal out_port_from_the_pio_overdrive_gain : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_overdrive_tone
                    signal out_port_from_the_pio_overdrive_tone : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_overdrive_volume
                    signal out_port_from_the_pio_overdrive_volume : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_tremolo_stereo_bypass
                    signal out_port_from_the_pio_tremolo_stereo_bypass : OUT STD_LOGIC;

                 -- the_pio_tremolo_stereo_depth
                    signal out_port_from_the_pio_tremolo_stereo_depth : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_pio_tremolo_stereo_mode
                    signal out_port_from_the_pio_tremolo_stereo_mode : OUT STD_LOGIC;

                 -- the_pio_tremolo_stereo_sweep_a
                    signal out_port_from_the_pio_tremolo_stereo_sweep_a : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_pio_tremolo_stereo_sweep_b
                    signal out_port_from_the_pio_tremolo_stereo_sweep_b : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_ps2
                    signal PS2_CLK_to_and_from_the_ps2 : INOUT STD_LOGIC;
                    signal PS2_DAT_to_and_from_the_ps2 : INOUT STD_LOGIC;

                 -- the_sdram
                    signal zs_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_cke_from_the_sdram : OUT STD_LOGIC;
                    signal zs_cs_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal zs_dqm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n_from_the_sdram : OUT STD_LOGIC;
                    signal zs_we_n_from_the_sdram : OUT STD_LOGIC;

                 -- the_sram
                    signal SRAM_ADDR_from_the_sram : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal SRAM_CE_N_from_the_sram : OUT STD_LOGIC;
                    signal SRAM_DQ_to_and_from_the_sram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal SRAM_LB_N_from_the_sram : OUT STD_LOGIC;
                    signal SRAM_OE_N_from_the_sram : OUT STD_LOGIC;
                    signal SRAM_UB_N_from_the_sram : OUT STD_LOGIC;
                    signal SRAM_WE_N_from_the_sram : OUT STD_LOGIC;

                 -- the_vga
                    signal VGA_BLANK_from_the_vga : OUT STD_LOGIC;
                    signal VGA_B_from_the_vga : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_G_from_the_vga : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_HS_from_the_vga : OUT STD_LOGIC;
                    signal VGA_R_from_the_vga : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal VGA_SYNC_from_the_vga : OUT STD_LOGIC;
                    signal VGA_VS_from_the_vga : OUT STD_LOGIC
                 );
end component VGAProc;

component sdram_test_component is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal zs_addr : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : IN STD_LOGIC;
                    signal zs_cke : IN STD_LOGIC;
                    signal zs_cs_n : IN STD_LOGIC;
                    signal zs_dqm : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_ras_n : IN STD_LOGIC;
                    signal zs_we_n : IN STD_LOGIC;

                 -- outputs:
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sdram_test_component;

                signal FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal FL_DQ_to_and_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 :  STD_LOGIC;
                signal I2C_SCLK_from_the_audio_and_video_config_0 :  STD_LOGIC;
                signal I2C_SDAT_to_and_from_the_audio_and_video_config_0 :  STD_LOGIC;
                signal PS2_CLK_to_and_from_the_ps2 :  STD_LOGIC;
                signal PS2_DAT_to_and_from_the_ps2 :  STD_LOGIC;
                signal SRAM_ADDR_from_the_sram :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal SRAM_CE_N_from_the_sram :  STD_LOGIC;
                signal SRAM_DQ_to_and_from_the_sram :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal SRAM_LB_N_from_the_sram :  STD_LOGIC;
                signal SRAM_OE_N_from_the_sram :  STD_LOGIC;
                signal SRAM_UB_N_from_the_sram :  STD_LOGIC;
                signal SRAM_WE_N_from_the_sram :  STD_LOGIC;
                signal VGA_BLANK_from_the_vga :  STD_LOGIC;
                signal VGA_B_from_the_vga :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal VGA_G_from_the_vga :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal VGA_HS_from_the_vga :  STD_LOGIC;
                signal VGA_R_from_the_vga :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal VGA_SYNC_from_the_vga :  STD_LOGIC;
                signal VGA_VS_from_the_vga :  STD_LOGIC;
                signal clk :  STD_LOGIC;
                signal clk_0 :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_estatus :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_multi_readra :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_readrb :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_status :  STD_LOGIC;
                signal cpu_custom_instruction_master_multi_writerc :  STD_LOGIC;
                signal delay_time_to_the_membuffer_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal in_port_to_the_pio_output_power_left :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal in_port_to_the_pio_output_power_right :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal out_port_from_the_pio_bitcrusher_bypass :  STD_LOGIC;
                signal out_port_from_the_pio_bitcrusher_crush :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal out_port_from_the_pio_bitcrusher_downsample :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_pio_bitcrusher_drywet :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_bitcrusher_flavor :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal out_port_from_the_pio_bitcrusher_tone :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_compressor_bypass :  STD_LOGIC;
                signal out_port_from_the_pio_compressor_gain :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_pio_compressor_treshold :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_delay_bypass :  STD_LOGIC;
                signal out_port_from_the_pio_delay_decay :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_pio_delay_length :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_master_volume :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_octaver_bypass :  STD_LOGIC;
                signal out_port_from_the_pio_octaver_dry_wet :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_overdrive_asymmetric :  STD_LOGIC;
                signal out_port_from_the_pio_overdrive_bypass :  STD_LOGIC;
                signal out_port_from_the_pio_overdrive_gain :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_overdrive_tone :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_overdrive_volume :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_tremolo_stereo_bypass :  STD_LOGIC;
                signal out_port_from_the_pio_tremolo_stereo_depth :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal out_port_from_the_pio_tremolo_stereo_mode :  STD_LOGIC;
                signal out_port_from_the_pio_tremolo_stereo_sweep_a :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal out_port_from_the_pio_tremolo_stereo_sweep_b :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal reset_n :  STD_LOGIC;
                signal sample_clk_to_the_membuffer_0 :  STD_LOGIC;
                signal sample_left_in_to_the_membuffer_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sample_left_out_from_the_membuffer_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sample_right_in_to_the_membuffer_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sample_right_out_from_the_membuffer_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal x_in_to_the_analyzer_input_left :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal x_in_to_the_analyzer_input_right :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal y_in_to_the_analyzer_input_left :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal y_in_to_the_analyzer_input_right :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal zs_addr_from_the_sdram :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal zs_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_cas_n_from_the_sdram :  STD_LOGIC;
                signal zs_cke_from_the_sdram :  STD_LOGIC;
                signal zs_cs_n_from_the_sdram :  STD_LOGIC;
                signal zs_dq_to_and_from_the_sdram :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal zs_dqm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_ras_n_from_the_sdram :  STD_LOGIC;
                signal zs_we_n_from_the_sdram :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : VGAProc
    port map(
      FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 => FL_ADDR_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 => FL_CE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_DQ_to_and_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 => FL_DQ_to_and_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 => FL_OE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 => FL_RST_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0 => FL_WE_N_from_the_Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0,
      I2C_SCLK_from_the_audio_and_video_config_0 => I2C_SCLK_from_the_audio_and_video_config_0,
      I2C_SDAT_to_and_from_the_audio_and_video_config_0 => I2C_SDAT_to_and_from_the_audio_and_video_config_0,
      PS2_CLK_to_and_from_the_ps2 => PS2_CLK_to_and_from_the_ps2,
      PS2_DAT_to_and_from_the_ps2 => PS2_DAT_to_and_from_the_ps2,
      SRAM_ADDR_from_the_sram => SRAM_ADDR_from_the_sram,
      SRAM_CE_N_from_the_sram => SRAM_CE_N_from_the_sram,
      SRAM_DQ_to_and_from_the_sram => SRAM_DQ_to_and_from_the_sram,
      SRAM_LB_N_from_the_sram => SRAM_LB_N_from_the_sram,
      SRAM_OE_N_from_the_sram => SRAM_OE_N_from_the_sram,
      SRAM_UB_N_from_the_sram => SRAM_UB_N_from_the_sram,
      SRAM_WE_N_from_the_sram => SRAM_WE_N_from_the_sram,
      VGA_BLANK_from_the_vga => VGA_BLANK_from_the_vga,
      VGA_B_from_the_vga => VGA_B_from_the_vga,
      VGA_G_from_the_vga => VGA_G_from_the_vga,
      VGA_HS_from_the_vga => VGA_HS_from_the_vga,
      VGA_R_from_the_vga => VGA_R_from_the_vga,
      VGA_SYNC_from_the_vga => VGA_SYNC_from_the_vga,
      VGA_VS_from_the_vga => VGA_VS_from_the_vga,
      out_port_from_the_pio_bitcrusher_bypass => out_port_from_the_pio_bitcrusher_bypass,
      out_port_from_the_pio_bitcrusher_crush => out_port_from_the_pio_bitcrusher_crush,
      out_port_from_the_pio_bitcrusher_downsample => out_port_from_the_pio_bitcrusher_downsample,
      out_port_from_the_pio_bitcrusher_drywet => out_port_from_the_pio_bitcrusher_drywet,
      out_port_from_the_pio_bitcrusher_flavor => out_port_from_the_pio_bitcrusher_flavor,
      out_port_from_the_pio_bitcrusher_tone => out_port_from_the_pio_bitcrusher_tone,
      out_port_from_the_pio_compressor_bypass => out_port_from_the_pio_compressor_bypass,
      out_port_from_the_pio_compressor_gain => out_port_from_the_pio_compressor_gain,
      out_port_from_the_pio_compressor_treshold => out_port_from_the_pio_compressor_treshold,
      out_port_from_the_pio_delay_bypass => out_port_from_the_pio_delay_bypass,
      out_port_from_the_pio_delay_decay => out_port_from_the_pio_delay_decay,
      out_port_from_the_pio_delay_length => out_port_from_the_pio_delay_length,
      out_port_from_the_pio_master_volume => out_port_from_the_pio_master_volume,
      out_port_from_the_pio_octaver_bypass => out_port_from_the_pio_octaver_bypass,
      out_port_from_the_pio_octaver_dry_wet => out_port_from_the_pio_octaver_dry_wet,
      out_port_from_the_pio_overdrive_asymmetric => out_port_from_the_pio_overdrive_asymmetric,
      out_port_from_the_pio_overdrive_bypass => out_port_from_the_pio_overdrive_bypass,
      out_port_from_the_pio_overdrive_gain => out_port_from_the_pio_overdrive_gain,
      out_port_from_the_pio_overdrive_tone => out_port_from_the_pio_overdrive_tone,
      out_port_from_the_pio_overdrive_volume => out_port_from_the_pio_overdrive_volume,
      out_port_from_the_pio_tremolo_stereo_bypass => out_port_from_the_pio_tremolo_stereo_bypass,
      out_port_from_the_pio_tremolo_stereo_depth => out_port_from_the_pio_tremolo_stereo_depth,
      out_port_from_the_pio_tremolo_stereo_mode => out_port_from_the_pio_tremolo_stereo_mode,
      out_port_from_the_pio_tremolo_stereo_sweep_a => out_port_from_the_pio_tremolo_stereo_sweep_a,
      out_port_from_the_pio_tremolo_stereo_sweep_b => out_port_from_the_pio_tremolo_stereo_sweep_b,
      sample_left_out_from_the_membuffer_0 => sample_left_out_from_the_membuffer_0,
      sample_right_out_from_the_membuffer_0 => sample_right_out_from_the_membuffer_0,
      zs_addr_from_the_sdram => zs_addr_from_the_sdram,
      zs_ba_from_the_sdram => zs_ba_from_the_sdram,
      zs_cas_n_from_the_sdram => zs_cas_n_from_the_sdram,
      zs_cke_from_the_sdram => zs_cke_from_the_sdram,
      zs_cs_n_from_the_sdram => zs_cs_n_from_the_sdram,
      zs_dq_to_and_from_the_sdram => zs_dq_to_and_from_the_sdram,
      zs_dqm_from_the_sdram => zs_dqm_from_the_sdram,
      zs_ras_n_from_the_sdram => zs_ras_n_from_the_sdram,
      zs_we_n_from_the_sdram => zs_we_n_from_the_sdram,
      clk_0 => clk_0,
      delay_time_to_the_membuffer_0 => delay_time_to_the_membuffer_0,
      in_port_to_the_pio_output_power_left => in_port_to_the_pio_output_power_left,
      in_port_to_the_pio_output_power_right => in_port_to_the_pio_output_power_right,
      reset_n => reset_n,
      sample_clk_to_the_membuffer_0 => sample_clk_to_the_membuffer_0,
      sample_left_in_to_the_membuffer_0 => sample_left_in_to_the_membuffer_0,
      sample_right_in_to_the_membuffer_0 => sample_right_in_to_the_membuffer_0,
      x_in_to_the_analyzer_input_left => x_in_to_the_analyzer_input_left,
      x_in_to_the_analyzer_input_right => x_in_to_the_analyzer_input_right,
      y_in_to_the_analyzer_input_left => y_in_to_the_analyzer_input_left,
      y_in_to_the_analyzer_input_right => y_in_to_the_analyzer_input_right
    );


  --the_sdram_test_component, which is an e_instance
  the_sdram_test_component : sdram_test_component
    port map(
      zs_dq => zs_dq_to_and_from_the_sdram,
      clk => clk_0,
      zs_addr => zs_addr_from_the_sdram,
      zs_ba => zs_ba_from_the_sdram,
      zs_cas_n => zs_cas_n_from_the_sdram,
      zs_cke => zs_cke_from_the_sdram,
      zs_cs_n => zs_cs_n_from_the_sdram,
      zs_dqm => zs_dqm_from_the_sdram,
      zs_ras_n => zs_ras_n_from_the_sdram,
      zs_we_n => zs_we_n_from_the_sdram
    );


  process
  begin
    clk_0 <= '0';
    loop
       wait for 10 ns;
       clk_0 <= not clk_0;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
