��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t����j�X�8����B��c�AϓT`���oj�~|��,�E����{���5�qȣ>�ub'�s!��^͌H>��50X$��J����4�ځeiz��eXIѝ]�\������L3�h��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HCZ�C�Ru�����[H��22P^��{������6�a�WN8�L�u�E�>F5��o{�R~�Y\m�Ȕ.��K�Q�ց2.����/8��cG��B�+�%Y栠��'ޭ�--j��7��ml.���~j�n����©�kh�ؐ��=?�^J.W�Ս�8�"n�B,�U��,�qQ�0��'vI�?�֐`6^�fv����x�Bڻ�.8��9X\�7������TиEm�;����ME`���͎�ݱ�tĳ�U�����Qw�_� �6Тj�&[+�{˲
���Vŋ3`��9b�ϡ<|�9 L�p����\�%p�+aNߎ��l�;�0�)��Q�؍a5O<�8k�P��gM5�5�+}���?�h��ᤊ7d?4��_ڼ������E)�N˴vU3#JR�'H�y�a�bC�y��r�%�|������D~e�P�����{�R�����φ1�V�$� �մď��6vU�An��&{\Z�/S�o�0���4x�.vtٟ��9�9�z#��q"�3���6ș�*t����K9HR0�䒨,�('�=1�3^��O�w����e�yH�6��xG�xm��:��_�mVSw��7�q�ke�;�f��^�����ް��>��f;Ʋ͜+G�V��ؼ�aL��6��i����q�������2b������ʦ�X��M%���$�Tc�<��m�2���p��
��l�0�cu^���ɬnDA��|g���C}��~��hĽ4hc�_��ޣd��*"��&����&8z'��𔯢���� Ư{LJ[��\I߼9�w�hz���p���W���"��6y�h�T'�w6�u� \�1/\SƬ�V7�y�Q=E.p���6�x�T#c��Y��O�<by�U4�׃Y7q�Ć*�NFp"1�hbUz��]	�+��MjGAQ��O~�|@���cv��a����^�ixŇ�:3� �3 �.�4J����V�K�h��[��O"�A�Y�
.G�R:����<%�ۋ�c�ľ�B�h��A���U =���ԟ����;Y�6uxZ�z�����5���;Q��T���q�v��H�hL5+̈́Hc_��%�:ڗd#4��Ir�~9
���&8{��#@�����V�	)V6}"�؞!��Q��/�ه��i;~O��΁=�Cgz�s�M��l���oO��MG�����N�i�)�&��UJ��_O���\�=�>�!��Cޗ�޲`sԋ���x�,���Z�;�h/���������d;�Ω"��p�^3J�SE�O�)�׸�a��p�*�잱A��)���TR�fj+�I����>@cT@�s_�:�{^���P)�/�sa^�a� �,4ϛ�8P�ۈ-=�_�x�R��׃IL\�o���.!0��9���ǞX��ހaVhАmTi���t�S�$h��:��:D�W�L?U6�����7�>�'�%8�s��łYF��.��	��ی�
��V�����Gf/v0�T8!ݓ��N��-�/�{���5��tLX2W�a*^
#[��EJ���M�Gy����ɔw���1��7a�v^y ��u!v��r�4��ғƟt�B��T!��L*���M���/�"F��HB^9xi�a���2Y���F�YOrD�ؿ2��6aCO�Z	�m��:;��91^U��4*�g�B��<w�OM�&�9\��� m���9��s-F�{�6��M��g�*ED��r�h�n�ϻ=�r�� �A�����.�Q(7�z^��1��u��`�v*�;�s7�W
��Һ�Oq����˃���_1�ǲT��t �~H@̨v���k�C��h�YD����;��{a��ӡ��*�#��Ǎ/�r��`I1�Нx����ʷf����Vހ��P��xSh�6~���n07��j�9G���tiJ�h�Č�}��_��"&Y.��1j����Y�|
�����*IY��m��(�/�l�G>�>�S��(���T�����~��.�O��9O�����2�0��S�ViQ"'D��d��6$��?��,�-j�8e�ԍ�T'Ӥ�Ie�Ͱ�Q V���Z�%��#i=V�/0����n�� ��~�s5~�!X�t�w���W�(���+�Z��d�Ph������m���E�K��6(��	�=z�j����W �h$�yGFQ�1&����x�qW׹]��,,��	?�`��.�p�V�گ,������ɘr�i�\aފ�j^�>����=4�����L@�J4����
��� yh�Ⱦ�~��6z�x}ʴ�it!`��x�
c�2��=�#�s����.U=��e�0�G���oG.6���
@�
ڣ.O^s�0�/.��w��ki�0B��˩-���&��i�:�CO�0�����#xA�8cF���LDe��1��ھ&WR4�^ `�᫏{;�^����.�OP�A�iF��b�m��/K�}}aA�m3Sc��WEz������j�.*���N�(j�.�#�c��)zJ��I�Q�Q\Nf��0�m�f�'���U�q���D�E+���]�L{p��-ʁU�s��w<n �U�^�e�ψ�����-��;"�!".��0^��g2ň�Ԕ��p��3��Pn�@��ǉ�)[��)��enT����#XY
-{'o"i���?���A��0~�5�����&�'-�v�Ft��4�SR*{O�+5$8b����]f�6�X�;�mF��A�����"/F
�]��K�9e;-�#�U'�5��qD���Ӂ^NZ�?��PP�x��>|0߆��Q�"�_:i�䢺��м��Y^tt��m�:�,���3@#��P�vR�A]��������M��E ��k�U��c#����H5]=/���ǻD�d/�ł<�*9��V��W����g�!ʗ��S՘����t��+}�R��l~�hrRf\H���,�j,�=*�AA��8d�`D���g���\�q0�k�ͧ�=y��g�4 �5 %��UC��;��9X9&����J�0aD��<p4�\����[s��:�1��j.*��E���.��!�eT_���Q�	�w��J�v�������Ħ�y��f�r�5�`k�+�����Q`[]�bK��UVK<'��Q:�F���|e"����x����t{P7k�9v.<����Ca0H�s]�:2f�:�_ؗQ�Sg��WL��\�_V❂Y���4%0}���7�i eG;� ��~����埁��Q	n�疞�'��S4���g:�˓`�܁\����|��0���~�/__�� �#VY'ȁ�c��l�/�De�3*h�lD�nZ�~�z����Sc4ĳ��5(X�m"9~+����wg9����|�O��D 	j{�����!� T��O�N���|G�%�\>���y`-�ܑ0�%�x��>m���o��O��-�h
t!l���wH����{���.�L�Ϟ�|�Qd�/�ڤ�,�������v�t8�s<�,��P-N�O�s��o5�+|C��ӫ�#����g�B��̙�]��4�8gK>��HW��!�)/�;�5����T�_q�a��/�Q*�3�E�`%�,0pԪet[����S�����I���4��I<2�H�[�fR�B�qMD�"Y�(r������`��p��{ �Ҽk���O�,��e8ԣ���!�;�V;�>�dW��k�˄�1��Q��nb�ip1�Hn�j���u#��E���w���V��*1�g�8��*�S5�t���2\�Yb,��J|��=,���B���4R,��iII���*�NTs ԡ�^R�Q���a��T�|�`b�y����,h=z4��\�#���ܨ���́P� �.݈��{���6aq�5o!$�*�B��ڥ��8 R[o���H����ɑ-��k���վc�v��N�&sM}�4E�>|jܥ��pԠ&�H���z̽�I��J�$��- <#5���u�c �����5��U�zf��e��?A����\e7K�:vԤ]GǭE6��^�V��SzQMFS� ����YI6=H��:�{|k�o����r	-�i,5�����/�5%�쑶�F�s$s���B-���,i�C�������<; ����۵�	x8x1�lF�:�����_Aҥj�;{�4z
���AQ�y2�7�:������޹��~'{	v�]N��O��/₵뀁p��;6�am���a�ZlZ�_˘�����̗�~�'�fENk���aNs���̅ �C4��8�vc���HX���4Ӷ�L���R���}�Q�D,��<@է���͙����fY����H�����E� ��Zk����q�F�árA�F�Y.	N_XM�H�&��Ƥ?,���K��e��{�m����~w	vaW�>1�{*a�%���)��} �0�t�r760.�VyT��Fa��<�������arzpS8v����׵�e�K���x��,a�r��:,r�=��⧫�!��v0:�l�Ԇ�&�v0�S �t�&����>y�͕�oJ���IQ�%��?rTao���8|��̻J�:l0�h�z��
�ﴉ>��XcI�>�����R�ym��Z�Ȝf�y�?�6v�d��x���ZU'�w���%G�C��r$%�u'�6�%���O���B"C��1���dD-���j�
�jDy�u�"{�x��h+�
qH-��u.t��ɒ�Ԍ8λf��]戽Qv�g+�tJQɣVI�_O�����.�޹�_W\t+#1ǂ����%\��A�1���2	�K^<=<�BG�$��9���E�;t'���{@��In������j_˘!zk}��l�c�R��1IDq���S�J ���"�8�"��	����ڭ$�T!W�RM�Jԏ׋�%W�4��y#�J2I_:�O7rݳ�Q�pn"R㝥�
i�����s�������˸=�V�f����&1�ƿ ��`�I�}�<�B�u[n�c���T�C�D���#��S��x��w-���$\�.�7���h2�$/qĲ�B���ϻS�U8�}��DKr�8�K��3��ZM�zZ$xg_�P�n}(��:< 96����F���H�U�6��O�N=���|�����$����
��b��|h�ɟ�d�c�܊�y0:��3��AFA������<e5�i�Н��,-�G��csd΋��e��<��.�\��c4�?3�b)欱.a�����xX�>��p>,-n����U����'�>���mn�&L
�Z�/r��5�U�7�� ��T�_45D�H� ��BJ� ՛h�"\zӂ���FPV�4_�i�q}~"g�N@��9:Ʃ���T���*O����֣>X��88�D��XB%�6�v^�I���a���C�p�;�h�	~����Vn��y�=z����|4���`� {v�O�o�ה�����ˌ�-�3���l4y��Տ��J�^��g�!�y��2%����*[���0b<��]�Z��'׬�'��;3��\�j��Ci?�&��kL��#�+�T
)P�n1�`<.kgmbxÃ�+����R�A�\z�jp$����>Fi����ԙK8�)� ���͋�u�#|RC��� )ӟIV�e�!0���#�|�H耚��C#4����N:���%t'��g�,���FA�wVM�dO?�5���4��)���$�On�~|�؀|������i���]1y���������6��5�;����k�/G�HG9�&��xa�z�tnX#(V��9��0��A��4��N�]`8�-�<�DX���C!h�����]�fy�����:݌��wS	��.R�6YU�iT*���^�E-��j�6yTT۳b��7�h�rd���&�&�G"���8c0�r��1C�s�{k(�.���l���t2F�_X�R���Rw�y�A�^G��F�jǨ��'�v�4K%� Z�w�`����)�x�^�������R6�k�'#�֝��������"!ӵi�U����+�o��|J鱗ƓJ�f{��g�*������9g�d������{�5i�A�I���Q�e��V�REq��&^|k}�f��v؂\n�3pc��'(Lxu�D M��L��.M���ع��m��˸m����#$Z5g C��䭙$�[�Vo	����w�R��L��'W��T���=�H���ڃC�K4��zwGZ�|SDv_��0�^��nU�_'yvc��2'I 6D���6<�]��Λ-�,�3���*�r����C` Gg���yF��s��n����ʦ��I"�Φ�U��|�?�+�ZZz-���W]8G�(�ڻ��Jo(����d3S��9� ���d>�-���-��:Z���Av�-eĵ��M�Y�!�9;<��sM4w���\�;
���~b�>�ܚ��+O\�K)�i����P�ՙ[T� <k!�s��O��."
�����sF:v�L>��^T�Sl Tgҭ��u`x���!����w��6TD2�:�ri4^;���L�{ -��-�?�?ϜO7t!쫋Ƹ�� ]�x������d��(F��:� 9���+�m}~��ԗ]�|�e�����׶R�p���^D�S r��e;�Y�ˠУ=x�97P�?��;G�`쨳�ʡQ%���N����.�[7��u2��g�Jf�܂�©�<k̆�X�j=B6��aR��ml�W�XrV)�툑j��	����AV5� ^�e���LTRHӠ�K�h���z8�5�]Q��WC��	���P{�.}մ��5O��X)vl�BBf�a�x�Ds�X�� r4n��<g_�S(\M�+�
�Z&���U0m6����O����U"�*;��A�+���6Ʊ'��ʏMmޥ�G =�4�>�j�,���Rķ2��P��h�[�'�5:��C+��Jʍo��
h��y)�6��s���VL���Z��r �	{�ϭ�/%�p�RDzx�V*qQ)�g_��?׀�I��_��(Kr��9w�s�}�~?��{���G'KR�m` ���2;�%/Gۧc��S1��i���8n�T���7��T��N<53֒���E�B��:�]8wp���i���3s����t'���WwG�,�^��T�R)�!�1����q.���T{��^�
�GDM�A~t��];e����	��n�զ8��6_��-��1��؎/T�� ����s�P�>0�!;����䠲�&�²t���.�L�y!�)��]b}�\���3�uR2�'-���NR�)\�m!i��| �S�
�-�.�����T��4y�`���k����!��^�K���H|@c�ĕ^_���LW�2/QtO��P&>�W�	T���ĵ<2�g}]��������������NcNE\���D���)7���Q���>)^�}}}�w�Y��s1��^�9�"]K�~Q/e]u!���ۑ5���\D���Ҹ+P��nƑ��O%�k�L����G�h� A�8ڰ�S�T��	d�������>�Y����_�3�~7~U�ɼE����n��=-:�d�8=�����]��M���J/>��x�dQÏ������i���s�k��](�U8�2�ii��)ʮ��$��9]�5}I�����q�e~��zr@���R�~���s�u� ��^mF�v�0h�:h�%,~`Ú�H�o�l���� _�w��.}��3j=���D	�d�� �OE�a���D�]"��5��/�	rw_���Pm<?��x�4.S"�p�e,c��7t*�9��ME���/nt���6�/��)����X����X��2�^:a�<C-a���:�Q�n7O���YNbv�����Khȋ��3ۡpbx����r֘n�e;������Y:�Y(�/�C���/shH�Ŧ�x(���o.�Gڛa���AXclX��O��L?,���jKaST�L��/�P�XGY�b<�W@�yE�&A�'�?��-�I+ۧS�_\"z��whm���|�6Wa":����L7�So����ɯ=A��^��f ��l���L3��N��K��`�V�� ���U+Q�����#U~����rf��U&4�� �t�g���]�4��u#?wV荇=��a�lzGC��e\��n_��@ښ'V�/r�1E�1����J�!�DAU;Պ�&Ⱥ�Q_���g�6 J|�H�6�9F�]q��4І��W�� t���w|���C�^�)���%�b���ɖ���� Q����׎c׿�-d�T%sq$ַ�?gPX�F�u:���Io;�	��x��^����o������G��3�1y'�}�`(914NT�NJ!_&��q��׸�Ws%]>:�ly���{����D��O�5�xs�Y��ª�1�"7��G�G��ԖF�e��	�gY�Q�ψ�r����KV��w��;���Y4a�V��0B@�+�C�0����k�ow�MX<oڬ1�і��� �F��{M���CD�"����4kS�Z�����H�+;�*tj3Lz�����Ե���] ,	�JN�;ȶ.�ZVL��]ؔv�<�8�Cwt�N�	����e����f[ܪ���XXV�>�@9��nBP�-n$��
��@���3�*9��a�$T�_
��8s۷��n�ESO�Z#$b�[F,R ����^y����}��@��'x�.����ԍ�
� C}e�F���*	v����x�-U!�^��j��N��pt�p�Ci��0d	�	m�� !�v�܋��#�2<.ѧ9���fCt��Q���i*�抒p�܆
�!�
LC8������QF�(�MK�-�g��t����M�җ�n�`Dj[�����N�Kz��J6ma��;������؟��d��)���w�L�h�z|�"�8s��j�'96��>�֘���9AӔ<`dS������&"��݌I[ɵ��� ����Y��q��Sx�(.]��k�}��O�*e����q�n��Vw�8zp��c���n!G�U�1���Q�.�)�/];R��J�V�ʒ�9-4�Hm�'�Qͽe���_4�Zx37�,���/;��~pg��m��^	��g������J�hE�}�F�;�o���>Q(��p�E[X{�p��_}��K{c�Q� �<�����/)���qt8�J4�'�����2������D#�.�D�E;�e	��W�f�O�`Q�"SZ�����N�t�p���Sm�a	�:=���Ty�<v�d�U��?e���#w��V:��]�i"�!~�*tIO�?Bb>	�8��D{^�H�š���+�<�Rdg!��~���*�Ʀ�7�Q며��fu�<����׽�7�`�?PbDS"�|-���n9L-V�s�����Ŧ-���
d�De��4ӎ��Z����������}��������:�N���j��zߑQ���y�bxF���.+^t�
�����2�]�Y��fI.?P�T�q`ͳ�� ��|(Dvt���oR�?�Y�TT�����H�I���QPk��߳���N��`�\�]�6�H�wL��D��'�+��s$]�ˋ�-`M�\B5H��~)w�S�7�џ	3rSuB��}ć&
\��K��Y�D���e��%5�t��ߏ������fc���%��)�ˎ�Sm��vQA�Y-��Oi�̗�۷��ȴzF��&Ra9�1?�50�ѸF���9s�:Ŷ�<wr �ݒ^�A�g� А=�h��Y��T��;J8������%3�e��?_�)i߭\3Bٵ
K���!��R�;�MW$�b�[#��6|iRQ�Z�玆b��׼�|\��;����G�����~���UBb �g�t�F��f��O�F ̴,*%���3���g����*��"@��VEF2�P1��m�(j��k�t��_f�&hMU��n\�����r��3�ږ�����:_�������2��`0Z�8%,��/�y��9�?�w�N
X)�5G�/3>�\]�0�Z��hb@�˹�WEDS@v�\��P_���L�a�B<��ĵZ�����F��Q��d3��u����7L��Uo��6 �3�����6�����S&l��^,��z���ƀ���WA�Iy��� ��9�}�[9Zui_C��5�Nd|�c���[K��0�b���4�kQ�iIh��ɑ*g�:2M	����vmZ�� ��}a^�/tjH�N��7�����I�&i4N,�j�[Ql:7E��VPˈ�~��$����s H���5}#DT$%�C�||(� �Mx�B��!�:�ͥ�FQ"uT��_�2�L|��w:a�ܚ���~0܂'�'`�x��!����R�	:�w4jn��㿔�đ�p{�����Dx9f��]�Lq��e�]�$qA斺Z�C�WүlZ)���|��%�*�P`��C�)��2y��f^c����yP�<��֏eJ|1-/����Η;��}����-di�[,��
�w?� �j���	I&�8�ȴ�̸��uP�Xk}}}7�~d�V����� �~��`:�8��Msb����Ӎ��ڐ3��n-�e{��3�)t#[����VX���]�41�{��F.!grgiX�zz���Rl��"�*Eڲm݆�і���'�&�ԃ�Ś$�)��ɯ ��_x�Q�
������j��*!���_����%�[gߊ�Z��(�`�<�jRR�k@}