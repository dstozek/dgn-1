��/  ?)��ݟJ�9�����Nm��X�[�`�������A-A}�٨�p�[̼_;R��RX��8Ftw0��1~���&��o)vB�������B�d\���VR����zCU��t���1"e�=+���?T��,Q�ދŸn6Cv��:�u�� v�c0�#x&U������+-�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HCZ�C�Ru�����[H��22P^��{������6�a�WN8�L�u�E�>F5��o{�R~�Y\m�Ȕ.��K�Q�ց2.����/8��cG��B�+�%Y栠��'ޭ�--j��7��ml.���~j�n����©�kh�ؐ��=?�^J.W�Ս�8�"n�B,�U��,�qQ�0��'vI�?�֐`6^�fv����x�Bڻ�.8��9X\�7������TиEm�;����ME`���͎�ݱ�tĳ�U�����Qw�_� �6Тj�&[+�{˲
���Vŋ3`��9b�ϡ<|�9 L�p����\�%p�+aNߎ��l�;�0�)��Q�؍a5O<�8k�P��gM5�5�+}���?�h��ᤊ7d?4��_ڼ������E)�N˴vU3#JR�'H�y�a�bC�y��r�%�|������D~e�P�����{�R�����φ1�V�$� �մď��6vU�An��&{\Z�/S�o�0���4x�.vtٟ��9�9�z#��q"�3���6ș�*t����K9HR0�䒨,�('�=1�3^��O�w����e�yH�6��xG�xm��:��_�mVSw��7�q�ke�;�f��^�����ް��>��f;Ʋ͜+G�V��ؼ�aL��6��i����q�������2b������ʦ�X��M%���$�Tc�<��m�2���p��
��l�0�cu^���ɬnDA��|g���C}��~��hĽ4hc�_��ޣd��*"��&����&8z'��𔯢���� Ư{LJ[��\I߼9�w�h]Gr4��5�������F8��.��?KpYF烨�ʴ.�3��E�ն'oo\\��������!*p�@��6h�������{� �v��5����S���a�Wp��k��fwTn���x �xm�o�ɯum���fc��f+��1�R����Lq�V��k	r&��MHY���s�wo�ssa��*�YT��ɮ���/���~�e�}�}��Db�1b	�A��3��}<9T��~�ծ�"�c����x^���,Zq1?�荦��-��ѽ�&�d�h��$�o�(����Z�N��j����;G��*��}�X�]���LI�)h�y�f�bV.�x���lO<����qj��%���ӕ�� ���Y�aT���y��^#ҧ2��
�؅rhR�y�M��_���Eap�kb�5��q�D���P���,�����p��ޢ��*��3��vA�F�3�1Û-��t$�����ߺ�{�ʲw�	LW���=�]̐���[	�]��-M�6y���o�"%�S@������HO�4>EW�!�N��t8�ku��b 7gt���!Z���n_V� �}�,+��A��7�bR���o� �^��Op~�EwUp{��>���S�е�ř��֧�G�0�/Lz�!����Ϲ�v�Z�d^SBŞ|7��]��!�yf>\�������� ���X�|'2x5v�C���|D`ͧ�޺��S|��.)(�+�vz����X[<��Ut)�d�G�`�f���n�T�G<Ǌ~�<Rb*�M��z�{�B�6g4CC�l������a�W�[e��:x�j�6W�O�i��C�[�X��~���o߳nD�}��`R�CCRFR�C��1�M5��$�l�(S��Q�\�m�a��Z�����8=K@T�r]����gA� 1U�W��� ��ɤ\��i��'c��U�m�����{��P��t
`3�<�[��6I�5NC�|d���P�8@7��0��Z�񦁏�,�Snr���~��������)���%Q�zTh'�s�f��ҚV���#��TzJX�]<��(�����"��1��N3&��f������i�O˗4Y�r_.S'��l7�*/a%d���m#8g6u�ILk�c �Mʿ?�ȊX歆%Wg�]��3�jY����,�"�ȑ�} PmCs�z|���Z�!G��O�ޠ�z]�* ύX�t�
�CP����̥������<��o�f�yS�f?����5e`��ֆL=�3d�Ǝ���W�[`��Gu٬l\����U���v��� 8�V��iPߗ}�r�-� �u�лS�<��<̕zמp��㣉)i�wa���ZVBh:'����~`O:�0��U�S:���Vuמq�g��W�n"�Y^����_�����W+����k&\C�����U�[����!0�UJ�~�h+�41�
��҈�s����m�c�܋{���I�C�P"{PLy�4������|WLig*�;|�@G�;�TMJ������`e^��˗�?��U�xz�Gj3�~ �g�Σ*�Pl���ս^� ��<'��׍N���O�%��g�����>�" s$�ᾦ����bYaŨ>^<�S��3yZ,Gd+-�I+��8�1�x:�fp�e�}�������$6+��4U�ќ�����^�7�����K�l"�b�|��K1�>�A�p���i? |Y���V}���gf���˿�\kX�ނ��/�����\RH;bn�E�����Q>WË=��jg]�� ݦ�b�UY��ӏ^X߷��Ŏj�\D�&�S5&�zc~S�W���I�+b��-��Sڣ�6�lά%���r{iD��W5g�#=K��!�h7�c�����_;5"����^���j��H>��gO[5���wd=V��Jm�̓�x����?"8�	��ҬҲ��_z4��ࡆ�<oU�{Z�@ ���\S�n��B��_��@*�0bgԗ>*r���+�O�X$4�9ZPg�\��
�$X�!TJ�L��l������[4�"G�3V�-�b�� }��yRW��M�������ҝ1���R�!�{�	����7�$,Y�"r	Gv���ཱ I5m(���tX��� ���T%	ף:�[o���)v̚
|���?��{H��7;W������+��q3��[K��r�EY6v-�����m���+�9�U:byl(&Ia�z��"ڮ��r�A�!LM��c����|/UI7�&4Aڋ�l0z��X�H@d���N�.q ߦ)�����;CI�V$���OA��` ��y�����@ߍͽ�<�����g�b���C��7Ӟ���&b�WF��J]=� {c��-�2��� �����W��V"�B�$6oi�l��3�g��.�a�0^JWs���$������)�^l!,�q�v�J����� <���<��T����שkGb鮿i9M�Tbh��F�qN��I S��Bj�V
!ڱP�W�	��Q`]vd�״S�6����JKfꭸ�~�扈L�|׉�{'&#�ԟ��[�I��`¬
�d����ov�&��Պ�;���J,.���������/��6"d��o������=&�G1�8+LV1�y%����)�V`��X�u��G����E����;gʛsQh��1���*8������$\���"ʻR��8a��N�a��h�rSEE��5+fGS�����4��70ڮ� [�J^�	op�M�B����c+u�+$[�m"�ȇ^�jЅ�%�{�V��b%)uh�B�5JT���
�3�P<.��%�Y�$���""}���o�� �~4h�cBڴ'7e����?a��w@��T9+Sݩ%�[e褊���(�F��� ��l��z%�: �a�����2���ܹ��IĈ@Q0�PN���`9Ɠ����N��)k�A��Y��n�`���dMZ�<�'�9r�mڞ���PJ�����7�����a�C�?'9�pi�y��p2�mŒ�̍��Ԡ�*!����.ǇEu�R�OBU�}��ѣ9Q��fE��{�*4�VBN1aEk1y%��"5T,�P�� ��0��Qq���y&�-R7��.��� s�D!/�M�x�˫֮�n�V,k	]�s���(+�p�᱒:���˶䔋���x�k�p%�h�Ab��;�#6�UOP�Q��t��ywT�5�m�0MT6�E,&H@z���*W/���l�e���VH�k��\�֚?H�r�?W���T�K�j������wd�iBo� h�ZW�`���qu���kF��߯S�w�Ħ¬y-�\���P�2a�$�0��A��tG�G�H��\}p�Tg�:Z[6S�<���U��9K,o�c�;�E3pg����cK�����%0����=���л��r��ܮ���)��#�}#M+sp��(�\�k1�\R���4�<�Ծ�7{��Y��* o�HA+C�O6�sQ��$���<^8'��ZZ�O��C�z"V;rr5���u��s�����j������.�+`u����������&��¢�4xuj���l
CH��#��K�c����?o��ś���i3׷�]��*��T@C����9���VêgػM�3/��i�V@�}�Y�ax�1q�Ho��Tz ;�X�C%W�e<��^��<�Ў��,e��V�Mx@R�����@ ��{8ލ6?��
�nd~f7��8��g�9ׇJ_Tʨ��N�x����{�شz��o�0	���1Y�9�7�R��q���u@�z�v�9����]v�&�e$��S���m���G��f<%W��8F����&+�V������r�cN�n�p� �M���	���Z���t����b�Tp���rRF)�hC���oϬ.3�u!�~�6y��1�`ɎB}����3��ֵ�~��q)N%�B5"K'��8���q���}�J��둊9M���j3�4Sls6'�ʳm�l�r��A6���S{Z���o�sUn���ˏ�#��P���%�V0�dl�Z�'�Pw]+\.Y��C�kA��"Xx����0�/�R�a�*��:�c��xIq;��9-\�+�j�C&�f�3x�z�����O��s���t@%��O���6�������L�CH�x�.�.T~�C=��.#Nt�4���q�@��ٺ򪊉��4�v���+��~�4;?�.��R�k�}�<K��㕦$K�{[9��(�:�Rt>/3���&���c򆈤���"�vLY��y���&rW��ݠ����p�./ ��@�Ҕ�5]c�/`�]-p�i.���J-p^'ߜ"�N�I��,UZ�2��0Q
p�Z���Կ���/XO��/��A��3����x؝HR�дr�V��.v9��]V,\�8rR�UC ��zǚ��:�'hz�QhɈ�WDPE#E�t�fv��3_�r/�^�)U��rg:�%��zb�6�|�c�j��x|��=��8J�8�e��&@\����%�S@3�SEÕ�N�=�\w<kY�&���_�}p��"�@�>�e�b��K~����1�#԰e�$���F��u(#]ޘC�����*[ͺ�Y��T���7��B *%]�5pɈ��&��^�2_¤Jn0l�Ű�!4���h����~S"��k�@��TȬVE@ؓx�c俟��x��[��n��j��C)^�ׂR���j��%��u�M<'�0PKk�����.� �c��ȡ�NP~�=s'Jx�V+�z?uչ*�u�g�P��M�N^�`L��b-��e+|Z%aU��w
07��
�j6pDw�v��<��3_���� r/+(�����(���7&�<��2����!��aN�l	9O�/9i�2��$>�����Ԓ��-�O:�e�P�����6@�#��t�o�3S �S�}�&�΃K�>�B�u_�E՗̗�� 3�i��6kB\�Lx>�!۬UL�r�O�׽v:G�K�ް�.��n}pe��l�år��dKcr���I�~f�Chδ��{���'u�|����p�=!�AS��~9~u9�	��J>"��&��"�ǭL�j
.���ӛ��w|�n'ND�b.��J���,��J�G�8a#H����j���
�����B�ZE.`|�\O�T(����W�֎��������Jz���ERE$����ݜ]*t�$ �*�Ȅ�(�WX4{!����»��h���]��sE+�Qj��C���~/�w��WΒ��[�u�J�\d�u��7��l�S�#'�M)�!޼Qr�Hnn0J0������H`븽p0��;&dtD��m���UC�xb�BUI]t������ �(#� ^�S�Ͷ:jݩ�x���	hÊ&ÌZ�]r��F�ʌ�D��LBVK{�׃�G]6�h$N�Jɗ;��p��-��6��K�v�3V�_�|D�IG����,��0���m;���{�
ޗ���n�w|�8w�na	7�=�Q���2���;��^�BӹWW`�Qnf���|@�z諾{�Y
ˁq�PQ�r��q�6%`ct߄�^Ե��^N�@�g��v������'/B�c�W���P��ײ���,l�=Ds��Er��FN�����w�R�g��+�i$�����G7���� $82��>j4��d�I��Δ|VC��d�KS`���ޚo>�m�+�3��I��7�V�S�	q�r�����k-6����KNm��a@Z�򙪾9U��ձ�o��:{Ҋ���r$Kng{^�/,�u�%Ea�w�D�ȗ���^J�Y��ӕ�����B�X�ח?�ql��Y�k�}�r\|�Ѣ���,��,K,��IQ-ឫ|����m�u4w� ����c��m���rm�v�i(�!��z.��[� /I�7�� �8�m�<F8��k.Y.s�	���u;A{"ݍ��� ���=���c����;���A6�dҠ��y�Z-@�)�H�((����׵k1�"�C�[��\a��'CW��-�s����߸ՌdP�3��4��H-�q�"�
��F��'�p�Du)��/H�[���-��)��!?sηA�L���]�O���Ƭ����PZ�#��	�<�K�t_�w��iq���+�1��O�sC(�6t���P!=��h��9�<k��`$כ<����'�x��rg�,��m�l�������b�2�p�*2X;�&���Ni������:�[O%�gJ��'N[�}�2SE��g1��Z�^>��Q��qd̽�L�>g�����\�^>KQ��u�B�-��BK��R��$���[/}.r��������<7�o�����?���^
��bP� ��|�qƦӣ�M�TNXA-����F4;�����&`�
�,�[x��f��|�z��'�?��"'$6z�� >]�2�٥̼�q���\�Yz�X���	I�bJc�E�$�u�ϿHّ�P��,g�B��x�\\���x��� �Ό��}���|+����;_Vh
<ʃa��2>݌�,Wh��%����̹v�鷼��߂�o�x/�26��E�d<s��B����[j���#��B��\�s#ն�=������.��G-1YF�������U��D ���BC�����v����kg�Im\BF���Ƞ�'���2g����2���>u7�iB�q�Iho�I�TZ� ��=�a�B���Hc�xqH�A@��ƍ6'��JL ��t��+��'��̄sڱ/��s7b0w3_�.��#K��c�GT� 9��k<.9��w�/}^�MX+4EvV.��ʆZ]<�ԏ��%��.)��\/�53��h~h��a?���\9n�R���J��L�+�Q��_4�A����-�N`6��R��v	�1�u��O ���������/��ݓ� F^|�w��[1�5��yb����7|�_#S��/�7B�ޭ]R�P��$�I
-��m�E���W���<�'�p���|5e�7)�N�7�~1��>�\ô��i�(�!����I�c��DS�,z�U D�u���6��2%k�V� mp�^q�]�a��c!��&�my�~*�amZ��������jl۪{I<���V� �̟������a��ȁ}�?c��4r�z��#������ŵ:����Q�Rr"�C��~�V�X��
��.�3�~k������Y%������R�߀��1�J�1�^{EY܄$@��{�3���aQ�n2�^�"�2�z�e�
њ_	&�T^�`�9�md���Prc�V�;�bv�I����[�6�\��uW|����#8.U��G�g)�Z]xHI�1��l�r�4�Ԃ?�M�0�q?? ��G�~Nㄭ?�� N8B���I�E���ͼ-�b/ω�����"M�+淸m#�L����Jy���B.n@�M�S*TGL�CPQ�o��h�]�S|,�E^�@��c��,�?�oӽ$�m���.���*a��I7��wG�RJ3�=�pw���6�*�n㆖Z�Y\c�t�	�}ժ�#K��� i$1����=�[D] j9y������Ŷ��f�l��|��:SU�=���A���T�T%���ڀ��k`D��k%�����`CRj��g���p�BF��V	��6�74��4<h|������}�^�PxR_Q��6yw�S�5�{~ҁ͍é�߮�t}�lW��C�}7��f����h���菰���8
�r�$k��!�\| �s�$�|��/��]���q�Uעu�����!]��sc(�ߔ��n�� "�(c��1X {�7�r0���}�Ӻ��S(�0���%�7[�{d�P�P���dZ�b4���y%$�v\q.�2O���:Иu �G����<��1���Ȃ���΅�4-�e��-�G�D�o^i���L*���~��:{��Q��2�5r[-Qݢ�P�H�*���]�!�WMZ˄�)D�$Q ���,��;��$��2��ej�
r�4�:���&e�bT��iF�^R\G�2�����&��(�%��C���'����4�8�&A�XΎ#�PGUv�b��P�wc^�?}�W V���=�mB�}�8D3<�1��������oM�!-g15�]w���Wj�og��,JT��J"T���}$j搩V�� ���� ��T��Z4�
g`��.yw{����_�]G�<R���N�&s\!�>n�)GT���r;l��C(�	�oǢB]�[�f6�����%[0� h\�<��;��Ћ�0BI+m�
m�[Xc��������Zj�̧$�C[Ԓ�@:��-Q�F# ��1�/�j�H??vQ|��`|5��G�����J����}�H�ͺ"А^�)�3Lf�64��r?i�&�l�U��YN��7����	K�]�����UWю:G(�h���ںxю��;&�F�9n �=�1<���X^ٖ�W7�೹�3xͬ���4aA7�;.�����s��i�U|���V�j��<�)?�Iث�W �_Z.At[�z=�b$3.�ȥ���]�54�#��qʽ�J5 h-�c�����<��~��s1�'�w� ��L_�&.�匇4���/`#',z���Y���\+��Z����`{�\�S���s��1�*�᭡���ժ
&�[�4z	�f�"E�kKo�3��$�[�s��=�$;�h��Q6���1�O�[�(Y��|�Vq���\�2�n�D�9���$�	5��u	
�:����r�}|�����)�&�fs�/�7�6�����$Yi�`bϘ���M��Y3lf�y��+�G�����
���D|�UE�7�2��l�[2}��B���kF�)X{�1�@����2��ߴ��Q�ъp4\�Y���e<���n-ci�����v�,����%��$�)6��c��wY�ʋ�O�>ᰘ�V$ǋ���w̚�7�zu t%�1�f��7�����.9�U=���t;���ˠ���ń������<�Ǉ�]'��U���m�ӏ��e>���8ǔHQ��r9����O���cD��[�1�,�챚�x���cyY���rLL����ށ�j������������y���7{'�^rM��1������Pkګ����#��;�C�|��h/�X�Qj���!]�т�F��^�	�I��׋��AE����1��QpU�vf�8�]:#LF��}L��߮)#�ͥ��|nM���ځ]Z��s�錴8�'��EW� ��,�0To���jV���>�,��qJ��	g�$6�K��'��R���R%�=j�Ɯ�'-��&ɍ,g���ц��3�&^�3���䎨���l�t3jn�|����[�w{2�`�8b~'
ʩj�*��������3�_>�;���<η�hF�mgn!��][6웲��}���]L�)��|��m]�a��cVO.�Ӟ����JxJˊc��Ċ�Y��\���f#�s�3� ����:�Z)1�0\����)I�]J�S\?�Ƿ����9eB�dw���pSׁ��؏���G'B�������b�p�+?!aS����@���5'	 �Ƥu�C��{���\NU����B�;}J�S�$'�mzQ�&B vjG��P u��� V�����©-xǝO.��=I�Pq+^��#@��@��y z��w����
���V�L:^@:�衫����@�ݺ7�A�,X�H��ƚ�;�6�3W� �����m̾��pV)��ҷ�T�w`��i�&����k�_��г�ۏ�4xZM�z9"1�HG��w)�Z쥅xl�Ao+w^1�:��)H�Ƕ��7���\�H(��P��h&ޡQ��.C>�{9�Jy�4�B����k!���Ɋ~#e�"αx�����JB�^ÞPf~Z�(�pw�2x���(t�z�{��B���z �����3X��A�qTV�8���D1Rs�(oח$f�U�kF�=$A��Z-}O�r��Ե̎r����
�)���ɷv�.���~�v�j���Cc��.La��wsuE#4NJ�����؂~!7װ���f�r���f:�Z����d�ժ�gqgx(��gG�!c��I��{�8�3�<6�Ǵ|��(:�-�A���@��(�{��#_ׯ��j�Z$��	G��5�eF�������6�3_3�>zS{(5�gY�H	�w1�f���sP��8z���&n��-K���|�h�	����K�<ӄ�Zq��űCܕ�~�{�Y�_���q�c;�;��93K;%���E=�ë�����Eq#v�z��Z�l�p`u���(��VH��|�VwF�����I�ڶ��D�\3�
���Gd����f�:꯫0vCUw\�{�����ʩ��3���잁h�����o< ���:���)mzW梧9ˬ0&�.�	`�5ڜ�v�ՙ����2v�K����Fb�>��"?K�A�&"ȳ��ԛ�i0����7�
��@�L�%�����PQx����G��?v��V�Fu�|�״[�0W}`��X��Ʈ�����kZ�7�M:�&R9��L~HQ��M��P���-C]E�{��V�i��>�Z�d~b�]�V�h�E�SEh)�S΋�a��=8��>ա/]�Xz���d/�a� &ꦖT��UO+nGG��}�M��\0�yI
�U�
�zY���~Fq�Oj]K�Ln5�O�WN:?gW�Bc�ΣDϔ�[Lz�|��b�b0zb��J*8^�b�.��Q?꾎�om�$���a@J,����tB;�ڈtHW��]���6d���ҋ�;h3�8v���)�ৼz^U|ޠ����\��cn[�kyv�C�����\��n��=�~i�H�6��4��a��,�V��k`ɶ�x>�/Ɛm�t�BN`��z��wE���<˭�AEڏ��"����MTxڙx��e\>���
���L2�9}�2|�]/�{��M���6��F����7�˅����G���q�h0�\�O\�.y��c�8?�m;�'H"�l�,J�p<�a>���Zd�-��+�O�7�F.�fQS�{M^t���^b^m�74p�#��D���-ș\��㯚�{�Ho� ��Aׁ�ۮ�,hL�l����lQ��ɩ0��3,)���w4�,]���K�&Ej��1��db/� $\liϙ�-ꊪx��̹%\��!0��i�!��^Z�2Q��\9X��q0Lw��e@z�3-;���jU�j�Z/f}��A牦�h	d�:\�x��-̂, }�`BB{���S"�>��h/��� ��T�)���D��$3G�IV���"�q[&:6���T׳v���tǵ|��J��A1�SB�r�S����g���	�a�0j�@.x��q����p�8��P�?�&��-Q#�A��ca=:����ز ����5Y�J��!��7���`k���o~Z�aU`;x���ƪ6������܆�b��<P�M?�5�L�e/o���B3���xi�N,��1�B�"����0�:��c��*�z�}�����La��2KB+N��7�~���'����w�_�|R�- �9Φ�+�U�%���3���$�L~�ń�iW���������=P���.��A�ϋ��d% �|�|����/8M�">�3=V	/��g`-
��ԩ�L�\,!)�2z�������	��ԏ�E�kR�s��c*󃜉�5��R�9y���R��arF�{Ʌ1��C�5\��Y=�f���1g�B�|��2��8���a)�s�l�3��Ub���aX�3	�&IZ`�6�kcP�4�&M��gF���d��:��`P�����s�B� T^��lU)}+�?���Y��餤�u�
�й�(��m���(Yn��kM,WӲ����4η�9 
$&>�<tnز�~Pp;��{��(�$Ŕ���j�W��	x���ʗ���4}�МƧ7��tUk�wW���}@�3\�n�=ɮ	��]����d��3/�@��	���'���]e'Y���h�i^c��r��gt=�暼��M�33G�)�-7�~��Q�A��Sɯy����rA ��4���E�r�����Y���H��J?� M1��J�>wz�k�n��~%�G�P��u_<r��O�!��[0�R�y��?�:�g]D�ww�F��l2;[5�&��ʒd{Q)A{����7�u���ox=+�Wd!�o��0d���SW��XϦ��Us�~~���R,�K�L�?���2�Xi�+ΘvQ�k����	�&M��CT#34�G���}�7Ś������*%i���\��
�ԋ��		4�-��5��H�	�Bz���`hs� �i�t�����3m�X��?a])Á#����b��y��+�B��wj��6���=���sӣ\����[i�FNK�����>��;�/��fI���Е�%����oپ͑����xg��+��;����yʾ����iO$;W���B���(�{a�wT|D�G��.��Ė��Q�U,?s�Y�h� 7��ݭ��ኯ���R��޳I'��`u��^p����#��y�vl�z�v"m9|��@8��	�U�k� yi��̸�A�\�@�漂9X�r�Qȡ4�BN9Hp)�J{���RV^���xw�T-���Ц�$MNG�C�#�]V�c�3{���dil@^�����(j��>��4'�镞��zJ��١љL��X�b'��0�B�4�M_�y��-��w���Z��<h<�u�XMq�Z�Nz�ɗ;e� 
1ΰj���' �)���'�v��r_�1�*�v�hQ�ߑ�9�.�����kH`T��?��t㭘�E��l���ټ�$��dÏ/ID��'V"ʿ�[�����!�3�%$Vh���9��/��I�CX�J��xܦ��ͱ}��ƳH�d��RF��h3&N�"*�n�$�/+'T��¼R�]!��7C핖�U���@c�d�3Z�aj�dK�͆W�O��3�G���tnXc�3�lG̮��I<�)1�
D&C�ّ?���OOt��5>f�e��XC�Y�/�-���,�i�@��t�r�۔�9S�x�3�� �d�#��W����c%��Uo��@H�t[�w�+�ǣ0Sɣ8���ɺe>��I���l,?���X��	^��Fqv\h���,Iߨ�u	fH~��f��1��@x��: 0��3��w\�I��V�%�cY�BV�ƨ�C�gp}�����7B^�;�I+9���6�#����.�Nl�؊f���,Z�6,�4��</�j8sӖ5�}�@���gv����;-��i�i�|Mt������i��p�y���� ř�u�.������B!k�?�����9�T�9�b�]Rꆄ<�{W���T�g�s )���$���3O�j��(pbs�ׇ���4�%��*�.}�m�|��_��'�p�J�LY�BN��'��g2�3� �U�xj�O��iĩD���Z^�3�
|�������G�ິ�g�;]�𞭕�3ݰX��,52�y����HZ��f�,��V��j�z�E��������͘�^���ֶ������~�\i;�b�C[g�.������g2�� B��{�e���l�)6Q����H�6�G���c����{�DK�/B�pa���"���+�k%���p�eퟕ��<���P ��D�~H�8&�?*s"
}�9�F-W�!�Į��B���+L�%d%�������Z^hc���d���f�U�w̺�#�YQ�����i���e҈ ����ܐ<�N�]����و���bǵ��/�XXo�oeh��o4vw]ڧ�U�vxFV���A;�����e���,����u�J��}J :��,�d�'�(]�Tc�r�����c�ڽϋHQZ�Y����o�>�V�Fh��aVl���{2�k�#���m뻂��۰��_�ls{��Z{#���.�"K�)kx&�{�\,{�
=(j_�����
�|���ʸ���Z�]7�1��޼,�x�=j����
��\�-(�t,�UӾ�4�q�ܞ;%�q�/(W6!�H�%�H�S�y�Al¹�oȗ�G�3�����U	�n�Ii�&S/�#$��7����w)��S��}�R����f�nx�S�bBv�c�T�vMoQ1�u�F�J|����<d�o��7�n����z���<Շ55<dJ~FY�PHc'Ī\��/��5 �R��y {FL����ڏ5�~�\mU��p�^���is�*P� ��. N@^�P�ggo/Y�O
o;����6
���6��!�j�����;�-�|buեW�6@*�'w�!�v�F`8�=��;}2T����T�� 5\��|dߨSdm[�g`�wM=�!WE�6�6vQ�̵a�mHY�=�w�|.T�Ĵ���U9Z6�. D6WiV�����Kp��=�Aы��`TdF�z�w�Ex��Ӡ��K*���|�ů޽!�<��Z�8�
� l�����zcf{LX��n�~Y�UJq���t����;��C�{m�/�7o��v�M/�99��W����o3�8�js���?�	&	{!����;�o�}��E�s\�>K��
�?:��@j��=����3�u�$��98�U��-`���a4�O�R�؏ZѓLg��ց俉�t�0�FDR��Ӹ�C���A{7�+�[;E�v�=� ���X�]r��/���E�}L�tx}	��zf�"Ҏrh���+�ȠM��/�5֩ߔ��re��p4 �e]l��4\+�"6����(���٤�;f�զf��ҹ.��x"Ӄ�m3/�v������E:�y�if��F7	j�F�d�"ʩ���hK�h�O�'��s�te~vn�}�_i�V�W��$X���,-A, �:���܂�:��@<Ā&�G��_j�37.sP�s��^{��0�' D�ih��3�c�	{�9�<�##�Q�9�*,O����G���0~�b;{]8h5_�gT��*k��6���#��c����PaN�R�nI4p��eVq8[�Ì�%^�r*�o�t}���X�up�>�GkH��"w��`�z�hh��������	�jG�"d)�HP�|2��߫�r�h4DʂbAd�;��S�W9A�⃥�)���� 'cm>������9Y$�RHS��Ը�Щa<��J�]w�9���fT��D*Lx5�F��[�Qr"�zCt��U;lq�l%R+^<\��@�?yq�K�|^�vN�뉇�[d�"���$ޑ��1RV���/�>}�V~���n]�>v��fs+�/<Brm��9}O��ێ����������_�����j� tz���G�ML����B�M&���}�\/��DΒL^���{]r�2�fR�F�{,P�z�w'0���\���i�|�)}o��Z��/��L;��4�S�7��C�-���KY��^p�H�6��J�*�J� b2��UW�HW��D��<n����9O��;`��Y�4r���Cx��9/���,���"�l�[MNs����l3�
d5�8ܳ:m�6�C��Wqb�H�+�3�aL���9����<�m7�/^׹9��7�1:
���_�u;�?I��&�����<���{�5��� Q�h��%�ʨ�w.��0'gLS6�ǅTX�cG$ܮ��ƶ��9�3�5�ar�}��(u��!�8���8���ƈ�<`�J�-�KV�)�!æ�j��h�