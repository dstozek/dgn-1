��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΡ��'�N$4b<9^���_.x.�S�}��_�wd�rV9Mz	kb�X]!��:J�#�7�{r��x���:ό���Ȱ�2y/r��m�\�R$�<�V�1Y ��\?;W^|�bAj������h�W<j4�U�e�c�ދ�c�k�1�xix�`J�_f�2�	�ӊ�Y�������-�#����R�9]#�G�QӠ��
�N�< ��/F�+*��?<��i�/����b���X*�ꂖ���c �c����Ҭ�rsoEAC�XZ�M[��������}21�N/'S�2��b� eM�x��44�hVk�
����*6	���ҡ���㛜�
��>�VCޗ��9@�ܴM~�����~���:�[>�!����W	)T�F³�.�sA�Z��R�a����F��S:YB0:�;��Ť��27Xaϙ*);���%r�(!d5cbj�!/Tל'�N�!�w5��f�_ࢇHڊ�U���W�q��)����b"���bM��T��m����7~�.�<!�o�0��`�ˎT�˼�c���&��;��Ў��<���ƞ��s��X�r�Y�����/a>��_�w����9i�#\����h�c0�b�\]Θ�%`�@] �:s���m�d��Z�s����F�f͜��p&GqC����ι�L|�P^L�&!Aw��x�9U\�+�f;�jI�(��� 4W9Lru?�F��'a������N~���B@M��bf�9I"ei�j�ySe��r�o��g��qP��&p��M�����(qK����4;B�y�>׮��f}T�"�|��f�
G��՗$��`p��Z.��T�F\4��hD���x��O������ū��D�'�N(cQR@M����饷���a&��3����~�~V]�"N����{O.���ת<}�pgU��Y[bЍϠ�g�_�̿��&�WA��܄�Rv���c� ���0t֛ӄ@��2ʅ1�AR�t�@�g�,dP�w-�"����5� ŷ�u ��ш�AF�|�:(�T�{�P/	��a����VJ몢n❬�_d�3� F��x��0�b3� r�q�]"If�Q�L��N��za��������x�E��yn���;�֙��P�� q�a��h�"oI�����>"4�e�4�)�+�{�ǉ3�\�<T_�D�&�5�����^����9i��{�"�f(Ub��`�{��`&��q�/���1%�IHzAUz����n��C�/8;��@8��x>�C��W��g��a2��%H�b븀�8lw����3k��EH�Vg��~�1��ٕҐԻCk9���_k�.J��I˼PCO��Ǥ�5���e�9ψ�Idw�)	xDA��T��*��\X_�^�2������0`,�?"?��'4�H!�L�<��㌹]�{AC��1�~�Uɾ�����\���~g��5����}g+�'��ru���~-�z�dQ�9�[����[��,�'M��tu�m��#n��<�$�oRB22m�c���L�3�j����;� d�	iY՜F���U�Ix�/$}��-ЈkX6l8��脪�=hD�����R��n�2E��G�'��'z�x-\�KRk���̥�	�i3y�~��e�'0M8Kځ�⹼������fT����Y���>�w)����Ŋ)��J@�w�Z�o��������GV8�f�e�,����n��"?��1؏0Q�|>G����)�q!��3����q�^Ɂ[w� �)6}}�_.����$W�D�P_���x]Րa���RNEU�`�@oc��P1�#�d��á짼 4 � ;����p�z�QV�#?�n?�~��s}�ѵz�N,hi�.(;lh���ΐ��fLYQ��Z¨�1�����,QjVb%����|Ke&(��� ��^��Ԇ����?���͸7d����-Ϸ(�M�a��PſR�.���R��ZI7@d7�R��;��Խ���ԝ�w;�X~xb�o,W�̱'���8���0QҏD� 6�$yA�g�ᢏ�y�I���r�;����e�h���G�X������d���pG@��m�9X	�o�Ōq7�ak�`l%r��&�|�,���6�,p��a��"h����z����-J���7/�W����$Ǎ��NQ��n�:�<���̈́aA�s�����6��������<U�D�|��_��從n�g��tA��H��-�!��b�=�
-�9��ϊ�����L�^.�~ߔI�����X�M���z�?XU��	��b@�`�k�<{���#��¶&煝��LR�h�n�\:�x-%��1�����b?�?!��1�i c=�'9{,�S��Op+��.��,&^/<��
r�dO)��>��cۇ���!~=���|�l�=�_�)��R��!���]F-�AE�|�rL��A3������2#3��w���eo3��J��@��D-6��cTNae��;���c>���)Ԯ�>���O��Ԇ�������!)��}	��&rJW�E;+F��%�KZ�CΔ'X4��M�dC��J�a+�1x?�(�-���"��g���G�\�>��Md)��Z/ӵ�P�ٽ��߽�r���5`�B���U�1-�a�1yճ�.t�y�X�|����@���,.!���$)#v[���n�R��f׍VR�8@�#��%"Χ�&���H�$�i.���|�`e-8>���'��#�����"��!Ov�[99�ʝ�U�aY!S�F���^U�}��U�'��7�xʔ?���'!)����m�b�|p�h�暻8D�����$��apx'9�z:�w���5�!����˦&���CI<|Y�8�z�ȩ�� �W5*���d���@˥�<-'_�d|V��d,��!�k����OJ!?ĨC��E�ZכD���?#Ê�;�C�5�e�dx]�qz]Ԫx�G�ѢqJ���vk*�̳�UذHv��d��ȧ�?��O���mv"C;�܍��}��{���f�X&�u���?�#�:�+��2f���^X]J�
3
3��~PgҢix՝Ҩ�I��W"�)^%aT�x�>e�OZ� �=���FPU�ř�0�^��������<h֮�c�l "�-�5�
�6�ґ�����C/��Ҏ+�+y��2�u�,��X��ğ"Az�b�l�� ������qS�9��n-O��P��$\�Mj:�Z���Υr.26+?eHčxYY�d�2h�����������a��Q}z5tfg���]��H��m����D��������@�xq�)�P�zT6bRv :s(�<l�r#��:]���݆(��9�Rz��O�v .�ɗ.a�㮋�c.^�{y�e��Ô_�/"C!���/��҄?���IpL����H���^�	���O"|�O)q���Ϙ��'���Ѿ���ǉ�Y�����O�7=����j�pl�V$KƦ�s�J�IT�N�3l�8�6�)X����e�����J� ��-��V`ek+��Ŧ�(8�dfmy����|������^��-���iD�R���e{ TM�j�M�>��/��*�`��:��>_�� r63��^��I��'�6�lHm(���݄ZSpc�K@�kN�94�s�5�b{�� �<�@��c*���h�C�P��>)?�F��%%~n�_e/'J^����>��� Qb��e���ԿI<Fϝ@�	1�v���XD�h/��#���xB�Z�\��D�{@#S��]�&v���!~��k^Jag({N$f����3�&(|�")H�1�l����3��ME�&�{��_�+��6���ݙ�A;��p�$y"o�E���x6a�3�+�84+N�3��кF��+(�f28,'6�7A��Ƕ�~�Ts\9�f]f+?�(��>���4B[XPx/��P�Y�p�������]�a�s��S����m���������J��� tAĲ�f%cN-^N(S1��j6.�aO�Q�`�b�LFg�55Y�K�bz�5"�&�TS��|�4p#\bfc����o8<�;�!eo��>�?���͏z�ArBSૐ��D�Q��v�X��,F��$�xU���T��@�v��J�P�)3і����!���eK�߭�M����-E� �n0W*&q��9��w���'�Y�b���.�",��E��wCjW����w�!�C��cʥ��o0����h��T���a%[�RL�of�n$�I�cXN�eU;� /����T��r����6\���;�=�/��@iOUI��R�nYW���"�=�s��sp"��e��>���3� C��]����`����Z��S�F�e�#+��7�%,���Q��u���cz�3��1zm�۪E}��U�k��b��ϥ!	d���\��n+F輰0�C߶<�kx{9z��Ynt#3c�"�D�oh�]p�w�!���{~��TC�8��i(�Ѡq^�U�Ep��r��j��C֖��i2�l/q�HK;�PC��H��6��\@t�p�nL�F`�-��H�붷z�&�2 :�0Ѡ:age}��%�h��Q����EÇJ�K錨�����4q��٦�?g�LU��x��^�� ��-������������Y,`*��Q��^�GMRGbE���3H2�X�h�%f��b���Y�J����� ;���{<�'��s�p!P��o7gVN��3��A@mzw`���1�uD���L,�����Ԗel��Ni�F�Q�z�n�և1��l����T�=�7�%� 3�G[XF�]�;~���|Y�uњӹ|+d���Bi��;֡6���������������k�'���o2���f�὜߸�Gm5�[�S�c���F�Z�~�n��^�$���&��UKKO�͵��5�֐�_-���J�����`�z��Ǉ��=���xϬX��h^2-�	D:9��w^�貕�/q�f�+<��[��c�,:6׎��8Q�d8z�1�j������>| �AԘAP?�龩 n��vC�� ��E����\n�V0�SD��}�[]F�?xZi]v�w��o�5�EE(B� �CL�SL7��I"���u�;[�.v��8��q4�)�K��ێ��>l���<�9���;��2ׇ�gE%���Õh<���`с[��r�W�xum�5�O��sqë�����TΚuE��D�։�hC�t��ӛ! �L
g(��_A%2�x��)�۰M��rk�U�o2;z6�5F�L�*Nd�dI��b,�>3_3��h�T2OW������n���:1� Zd-O7�|��JΧ�5D>�����c�ވ
��8�,��+�����EQ��Q�q��9�OT�^0k�i�P�mK�v�)j�6^�~ǆ`vVT8��V���j�m̀B*�A�yq�)Qբ	��>�ޱ����2�,&3��P05d��UpY�M^��D���ۯH����ణ�uvj'%ǀ���_J��í��76a�N`]禸ʿ}�e�[�`nR�~��͠+~�W����´�S�s��Wx%�up����C�l�C�.Y�ʚ��w��(O�"�rj�?K\
\�W!���������kgYV0�E�ϣ9���'_�������/��b{?Q��ܧKVo�H%���uD��5��Ч{� ~d���K«<��w���@'*��5�-b�(_Ȫ�]߼~浖�o�6 U�������?��>�裆�yg��Gn4<��j�?��A��FY�>�{�-9�	�v�}u�Q�X�V���bu����k7>�1<����X-���x
�u$�C���j��t)q={��.�L�9%
��*#��:j1gl�	�pA(��d�������G4�!�$M��Vv}� ��v��/��v��r�)J�K�FD�y���u̱��x��ȉŐH�t�!k��I���|�
�i|0`���!������C��ȕ;��[��U���B�(i@$?|]�A{���9��/N�I��PU��E�OD 4+KԬ�"��+�c���+�8|��ȆX�8-����A�P�z��n��h���7�Pj��Ԧy�'��@��	yi�����;�����y�|�Cg��K��|���8f�����AYL�6��Ygk׊�g9����t�=�6)އa"6��Y��I�q'�8�L��+Ejɾ�'&�tѝ� �υ��`���l�V�8ݬt�{�<�@k�u �"nN����6G
�Ҩ� ���XbA�ꘔ�Z��]�sNSh1QW���л��>�����w�[^xD��R`a� 	!�����;KD����ØC׷�7��a��N��qu�?#>��_����SJ�u�T�Ds�)zCt��?v;��?�����j8{�L-�6/����"M�W�����&T��VqM�_�ǭ<̀�]�ݢl���~}�>��K��C�VMԻW}��>N2��2��X9	��P����,; {�	:x`���S��o
	S��ƞK�?�q�+1{�('�H�%������$uQQ&G���fq��`I��-_ileM�&���v��&*]*�i�!���[� U�Xv��86�:{8������5�k"�

ML�O��6����Փ"!��"%^�V���-^m��d��c�?	��?Տ1�� Ou�:�"��R�&l��%ne�~�����Θ.��̤�Z���9euI��B�=�1�dR;���%�|)�x�Y0�Vے�\T���Z��yܧ5���th��`.���x�+�qU��e���Bi��!R��YtԳ�ե��	�d�����Qr�YH8a�Q�F�ԥ��vΰj���yؼMn��v�^�{���MM}�(��F(�x���m�"?��Qt:VuXxݛ�RȾ%��XV���W�^�`!�q��l\ݜ�%x�N���&T��H�''�ݘ\K��@<���6����+�D��1H�����th�dŻ�t#�)�5�]���M�F�.��������.�l�;Qz~R3x�0�3��:o�k�f���X��G2@,���V��~������e�] 4�%OOq§>p�oZ}EPT���M^�5�ʲ�=G�"�26&�+o�7D�Ed�X5���!ɰ�Z�&��`��]iZ�|T��p��Qˁu4oa�`V�!-(��P������z����!1O�����z��A&�I����t��[�h<��ߑ46��+YR4%�Y������!��{�N��'\���n��
�D�`��I[V���	p~+��ײR���0Ϋ��<�;,�]�^�_6��ULa_s����wy�(_n2,�v�_�u�R��F�˨�`�,1�tg8�);�#�Z~4H�A̟��J${]A}�������irJ��w���"���@��&^Y��U��B'��H��t����I2��w���6Y����8��?�رZ��,:���p�0�~�'���C����g�S꬙OF��jeA9���8Nf�]]k��]�3j��g��s�{�
�X�=e*��*Ocr�K�T��^�`I����d���֓������8��<�&�ƍ�eg�|�sV�J�v��,]M�AM���D��ݠ�F�}j8��2��>��%�.�X��M��!뎃�����}��IPa�s&��<�{�y���/v��gr�L9ӈDĐ]��r�*��%-��Ξ�[���q��s=,��
�<C?4��U���HW��VZX1}Z������� �K�Kv	����BEA2͡t�V�S��)��0��S~��ǝ��[/Eᎆ�4;�=?I��u���S6T~�I��/�����iO��k��s��,i_Dﴝ�$_��P �1�����d�� ~r�F����C8�`x�)���<�Qi���D�m�!�<7yŸJ�����ڱo���n����
u�)��,��x�L8��L�GG�Ɠ��'8oti�1�t5�(͆Y]t�I:���,C:-9s���Bw�'b�S���.���R4zȩ�~a�P�}��	}-{�O�Kz�T<#h���Kq[jj�$��g(��u�4���v(\��|!��*h DX7��*�Ir�C!�W����V��Ύp��F��b����n�g���җu�$i��Bh�P�C:����=��2v�6,+��Y��Ɩ�R��tk�@o����`9R��_A�J�����O���*��ç,������ٮ����ë�x�j��g�:k�����֐�s?�)+�}&7��7�)ZPF'��ȯ�;�[�LZI��i��j=��,��]�o�9������j_4T)y���g�
�@���zd'أ���lhy�xo?_7:�_�ko�vZyk���_Vi���l�����h�sG�B��^E�&� ?
�:M:����Ʌ����mU;� <�8D�qq{��ҳ����iU�X�g,�L{u<�ji�������chuN�p>u��Wȅ�9�D�H��p�����0����ƅ`�=<�Gy<�
>�Aj���T�g�<f6-����$iAPvr�wс&�� vB@��s�|��d�g'7���5 �b�HC'�Ӿ�ێK@xR�h�+7����F���ܲu|~����l7�\=��#zp�5�0��z�;f��/S��5���ɨk�mWP�Y��˜����ͥ 
��/̤����k�Ȭ���r6��=Ln_�I��iI�׿��V��Q�O֐
Ѱ��|
�}�������7�GJ��|��ҶN�5$>p�<.#���W+G�^�\��.�v�P9#N!"Z
0�nl}""���M���Y��D
�MU ����(h`��6�./+��:��bX���g��d��H^uף��T9�i��4�R9�Y�	-�s�8��z�z�����C�|�����¥()�����'� osm!����%�̕[�U�?�']���W|�c�������Ϣ��j�D��,V�2�^���h!8I8��'h ��}"Q#�y�׼oS�/o-Z�{Ϡb�V ˟v�jL]�؂���o�G�ڵí����a�����	����Dh��K?̙ue��uq�Qd�%V�+E����kD�q)�n�����ٴ����1��cg�.��&�.(_��L
��(��(s-+z&��Yc���-�}��
�.77��#�p�ڡ��2�܅vGw�u�xGAw��S{v�J�j�;_4��p&�Ѓ)�K���˖�'>��b<�8
	t�i�
'fI��(���.�_E��㷧��lj�������,V%w+���I=m1Aw��zk�3����b�w���y�".))��9� ����O������rY>���2T`��K�X����+�Z�ZGH�l�qy�d�Q����?��W�y�wl'��v�M*��7�Ó!;�G.ѻ�[����c����D.>��	?��9M��	���#m��(N;3R
����z�������ߣ�J�4��P/�$�.�
�Ρ7e��y�gj/C�"t���ݣZ�Bj�J���i�J;8|�Ř�:HW\�s-��UE��yzڦ�D�c�6�[�h
	`����Gc��g%{��D@��ָS	��)�X����/=�`I���@�@Ma���h��=�-x�A�-~�q(�����,h:�QD�e�Sh?TnC���[�v��ta���\:�����Z
A��|�M[,�Z�6l�0�]�����|��ۖq9w����:��Q�m��D�d��:���>�  ��(��*^�d�����ԧ�ׄ"��87�:v 0d�s�m�y�Ĝ��7!���u���Z���\M���}߃8�rnf��}�9��f�On�锽6@V��x
D���H�K>#�l"pI
�&�e����Okeطkm><u�-��Wű�i��Kr9��DW.+��H���a�æ���1Ÿ۝b[�Ls��aA�R�t^����ؔ��D	���w�OJI,*V��
�X�uU[Z�W>��0R�<&���@M>ªg�>�p&�?�K�~���С^;/�#���0��+���N��ϩ�"�v'��>�y��Zէ�ل�5�yϟ�s�m����(����f��pAf�a�Z\,/X��8!�[ <DF�`X�6w�	
�-�I�+� _�JB��������3���(�kj�����$ėIl�hj-]�����ߊ�[�C��&o�Z�g�p"�v �61.�4�\n�V�J ���xa�M?�w���Vl�Q�b�'��t`gAMb��1S��;�!�v�w�������:�؜7�rh�B:Vʏ��W�49	��?�p;������t�Y�gB$��X��3P�ULr��9-�W�B�V��L��Ӷ���*����l�|g�"�.-�4��`-��mQY�OB#}p�r�uwF�g|��<ŤF�TA	�X���i���2D���U���`K��mKe��#��@L�>�LtW��5��GB�;y��qU!3�� <��@\v�"���E�8H>�L�$������?���'=�ل�y��Vj9��2��{���0���ٍ N�B1e2Q�a*{�ukHۨ�[�;Y��?7��p.�$ (/|���v��kf7�-���CWqkx69%L5+�"�����}B���O�מ���u����A��h��>�t��ע:��i�ȁ#�N�.c3����p(g����n:$�����s�%/�<z�t�Ӛ�!�)[s�+ .�Hu� $���C1�\�6���<$� \^g������<�*c�`��|�P+�؝�`ό����������f��5�'��c��g���<�MDF��3��qH�'O(I�G%0�q�k~��C�b$5|�m������PF��,F+.U�.��SC[�v�ʺm(o�ъ�oOZ�BPX�Cw�q�~U${𛒠�v������Re
��i)�T���	J�\����y��q�]���D;��y�������9"�:)=j��*S��:���E1Ӻ� �S7�ղ�(3ӾgdΎ���P�qy=��t8�^f��ZLK�|5���E*y�T=&�<���0�m�x�S�R�H7�4���i�^�4�y`���O��Q�7Z�L��y�(�^ G�F��>Lj�~�HPь5����������b'��pTmFTo�~�7���w�W�d��V�\ ��}95|R����qӪ��i����ƀOO�����\ͳ��}�Ԑ�,��E�ը�%��B3w�,�t��^�Rv��^Z��'���̛�&kfVs��	�j��׫E�"���n�����``M3����Ĝ���\w��t,��U9�K������w_(90U&��Q�x ox�q��{!1v��nx ��بs���)w�Vl��/�c��C�����v%�����NS�e�%w��� I�M�R���B�څ�i@�4�1�P����3(.^n���eL�@�5#M0�/E7���v�f�*F'sb���	rH�p��R��\߼Q��e{�)gE�ㅲjB�H�Cgky0z��]��:��� �=@�?�Ey�ztO0��|m"N/#h�Bq���A�ݽ!X���۰�D7��)Բw�S=�#n������x��3+{��;D��N����f�1��4;Q��w<7ؔ�R�n�;����Ǫ���U���� ��� 0�Y����m����U� fp;�y~hi��.��׍Q�����B�O͢Cn��F�Q�>=6�@�,�E½�^ȭ��l+�XC������}O��ʄ��QAy['�f���3�.�nq0a֜]V)�j�?69
�s���K:�o��cq<r��d�f!#t���
{r�k��` �D%B��F���!i��j�c�(�=���U�ޘ�.Hi+���5�N~��ë�Y�9 P�%n����P�)?mG����524��}7���/����]ްxנ�fY��ž��o3ms�<.hQW���(���Y���Y=�r�D���C��Y�=7���f�B0ގ5rJ$�����vR����@�fuc	-@�Ͳ��^66��8��z{ ;�@�(�sr<��L�Ph����ᑡ}�x�L�[��:�x�cT��.��~�����x�������|�맚Fk����
�ζn�Ɠ��?�O�����R4��X7��{j��<-�1kD�ʫ�*ԕC�\�	ǝ�_��������7��Q;b:�-A�w������O���d�u�5�7�<OǊ��5ʍ����H������%�=�R��ޑdI�k�`d-jz��˂�ݾD�7&v�o��G;|3sj���(���%�Lan�r{V�*k�q	r�o�S[J���K���̗��t�.�q�;��aӍB��#96���A4`�fI���*��Q���d�Z$��f0�n�S&���3�&]��bl�)`Vְ��Yl������/�I9�?͢dk��|W�,u?�IH�U3r�,��#׳�#�����}[吃���5/n������~Q�k��z�ZBC�`-	��A#`o$Z�Vb���
��׮-?��p�d��u9ߞ�zM7�\$~ ?W\�H���ۤ0����Z\�$���l�I3�k��5��v�ʄ,5�c>ըNn�>Ӂ���K�1m��]XӶD��<$*m�;O1G�v��8
t���Vq�p�+3�,Z$�N�tPx��.܏&)��hmn���
U�+�Tb0�g�|�·�5����{^��f�#����p+k>�FyjP��ѿ���%�S�@c<R�B�����L�z �����Y�f��������6��ᅠB0C#A/��u��f3v`�`bFM�Xt���@,5d�M��>���Aw��\n�p<v1r��<$��QH��[3	��
O{j�1a��1��@Gdl�jι�
�Z�I�ou3�j�2uqܙg�l��f(��~������eZN�	���O
/'[w)⽾dE]oU�7���4E�c�{~���
�q@-�z�"I1�@��|H{�.3J	c��+)�S67|L��|�rW�@�^%��Yl� �|It����8��Ǡ{��vl���K|�'�	��Dc�r��T��'"�+&_��z+�5�ze�n_	����c�V��.G�O�����v{jl/��1�����a��sB��~��H����c��5ު�r`�t�ِ?1��Vap�H�?d�����g���Ȼ�.
�̾��B�^�HB�M��g���kð���
��3nE�H�t���2uX]��wO�HaU����zZew�֚H�%��6�ړ��݆Kʊ�qG��?	��\�i��b��	
�9�\������_���u�}`�KF@q=�T�o���G"aI~l�c�.�9��!�kr���ʤ�E����]���-�*%U<v����f{��g�c|�hB��>�.x�yX��/�/.����j���`=`Z�k��빉g���'UBA�z������JqܙU4(�e��YOjs�����\Yh$ <3���L���.���{��U*��`�<O�YyYu����
�t����c��i����|^�N��R����5b�!@��3���@q���w�>�R��!;a6Mv�IQ�Oe�B�pʣȊ���s`�G-4�B�|G���ǨOyw��&Q�͖�ctjb�T��)9�E������:�5��ġ7=>�H8)S1.���Jp�Z$W(�9��y�LY�7I��p�N�]Ѵ���v��k�c��c��r�WN�6������5�u�g�	�������D<)�k�ksN_���#>����3���rqz��B\v<)]CPRna!������[@�UY5x>�D�b<0da+x�		;�ԥ����I�ք�Vs~T	�oO˥�/q�-:|.*��0��<����P�i9�An�|�֣�A*HZ�	����#���T�t
��D��Re�H�n��Ga,�? J�W��9s�5;(m&��wË�4�|Q�],�i�`�fk��|��JJg�f.��0�5���ثT�LĠ��r�����z�k�=���k���s��x9����wz0_O�9���O�ԅ<��ҧ�~��лm����O��˷^�n�R����?���9��=��t�s��
��ԇR��>�X��������D6�}j��V��Ƽf���;��?DI&yW�!zF�y�4ih����-���d��/4>������'Zk *�k��=])��`��e?C�X�T��ǉj��_�Ȗ�� a���	�s�#�@A�׫��;�ȃ����Q�=� �.�+�N%������ًP��Q�I�Q~��.��E�a�A���e�&�����N�=�	r�"��G��*^�k;�bmZ{,��B "l�=�]	pSppt�Ov�!><�a=�IO��P�$�Xf2ܦ�8}�nK�˩J����ޠ�#��RULn�6#*���̓�m������vFd̛�V�5(�V��ҵ����^m}����@�?���K4����vP�wO�׶�y�.�]��)~��ұ�)�P���:�5D����m.�[a<�\���4��E��}�,Suo�^�s������:���5#w-�	c����s��)�`�!�q�w����6�Q�^�S"c�������8h9��^?�}w�gE_�`�H�97�MG(��HE��p�Zi��� �,"�_*<@8�G�5@k!���yh~���Π���4ű<��'1j�O톗 t$����ZQ��\s��U�XQ����P$�����&��S �O4.&E�dJ�;�I�3&	��#/��F=�R���*{\x�oŠ�nh��3�+��unj[���&s������}�u�!��VM͹��l����L�B�:�0h�'���e#�[R]��R2�|d�jX�}h�v��(�A��=l�>౛)7�~�Y��m�ee���H��g{��߀uҤJH'�����X�i�2�sc�`ox��0ܧ��mK0�`O�ȕi�8�[	��P���,�2�#��yD� �k�V���1������A��yfu���k�6�w�&�����>kb�߻F��_@A�x����`q��1_w�����Ss)u�٘�����	��c�� ����ֆ�g�ATN������q�5)��hs\� �[@�cB< �!�����R,-~߻�FH|�q�V��@��80i|�6���>
��*R��b�=P����%3J�x$�iX��K�j��	x��ܚ4/{�2�n�7-D���lA$D��>Q�f�X�k��#V����D���(��$�A�a`/�%�z����-�$����J�UK)*$aM[K�K�S>uj�@�R�݄:��rI���Z|
n�,��`_9�UTc�Z��;��X}W8��5/����H(� Ԏ�l��m�-W�z}s�Nv�FT\��i�E���:��A�_嵄��
�$C6J��u���'�*޴��F1n6Q�3 ڥCP�{^g�#8�ʌ���V�}�SJA��sa{�'���>)�����L ��d���Ĭ��]1��Ǻ�{�R?�J<����K`P4�5�Ȉ���]�q��пr�]��A+� ����?e���>���{�$��NO	endf�f��\�����3�	�a/N�8<�ИNj�Ϣ��N��r�Ҽ=�D��/2؊j�]k�C&�ȵ�j���0���ڄ�g���┚��5��95����U�K���.�kdȪ����4��`!m5#��S1``������7��([�P,(����d�WدO�tV��&��H�B�)r��@�c��Y↷��ԜP�;Q[�����2�s`L`��"�_�a_@l �1B�K��rÿ�#�E}��o���INK�<��z�M��y�,n_ ���u$#^��{i�g�#8����Mg2W�(��iߤ�`w;s�4��ebB�At�wT�%W�%�	%ʼr�p�O�~�6�=���j�M9X�=y��jWQ�0?�p0��h#��ɳ��J�����f�s�TP��ԫ)t��ػ:����������
��Ae"����'�c�6zGyUq��g�4Oڡ�o���2����Pq���u���e����!;���o�Ho] � 9�_Z)
,+�顒[��n�
��~��uR��Ƞn#�l���o�	��4�~����.���CӃȎ�6�3+_��A8�{�0���f���ە�R�f���H/I �?V�%rtuS��?�Y�fC�P����||[n�!����b�9n���p?i1bz��<t�k��Z b��	% �{-��W}ފ���a�R���(L+�꼄����6��U���Q�q�+"1�U1L��6Z,I9���"����-L�@���n)��rE�WDh�e���a<�<%���j쉌����LOm�}h����G(ծ?��Lm������5jJg`�%�l:(H٩q6�(%r8�C�d&�<�d$��V�(���a�Ń�O�9�1뢡���d�Qׇ�De�_� <.q* U��՗�n�����$3�C�w���#"C���SA�xbO����`ۻ��ˬp�ě��oX�$����p���D$q�����L�1�V��H-΁�@��p�FG�=��q� ͝�\+Ap-�~W⻔
6͢ם��x�s�@�ko�5�%>/���-yh3v�/�w()�����Ȉ��f06{H��+�"y��d�8w��(
�/C
m#��^��7��@7�5,hGX]�ۢ
1|2Y|�͞-:�����#��b���a�n�o�/8�:���̓�ގi4o�ce-P{�P��f��Fv�7�Pt?+#.��?�R)�5�		��u���V�d:�zb0�e̓F�@(:oE�b�"��G3��
aw:���b��=k:l�n�9ߞ� �{�e��Y:ޕ�S��NT���hPD�u�Enc�aр<ef�D��!������<=w�3O�4�@�g0��=�1�ۂ��B'��^%�!C}����U>y��r���t6���+���l�6�"�Y0'�kL<��wJV �`T~��v��^��jľ�8�����s8�T������*队���)(�"CF�˅奠"ӸHE���o,�[��ȟ�ce8[����6|I{�@���Lmr?�L_��~T�# �e���)���|��ILFV����e\R�#�+r����(��P�����.�|G��|��j���C����.�_-E�Wax�I���Z�i���ۊ��Rc������P�n�3ޝC�|t[��DV�V�/M�bfw�l k}�㾅@{��;n����ʆ��{�U�HK�J��+3<H�	h�C;���
sǌִ�����5�����z���^C�#�o[��#����;��fFO�$m4��s��T՛M�N���'�4J�D�<�Ft�����(�v� 2��9[�+Gt��7]V�yq���o�D0��I&�Q�K�s�Os���.��:��e��K��I���A�1�X1��0��+O�H�� �UԏwM�/7^�^�@�\9�(��\�[�
,,(od��'�%0��7��zE����%~����8GtaԮ�2��=6G,�bBq.+�	��,�aϫoх�80�\$2���|�74S#[�E�G��ګ�#��s$�&�(G�-��8�Hǵ�|;^ЫO��g#BlK��A�����h��.h�� �_�d �r��sS��Z=�H���$�t�\f�j�ȇJ�,s�T�p��ٰ���j�GzP� ���N}����qh�%�ڈ��qg��	�?��S۬R�������,�~�'7��@V�Ɓ!9����p�O�oK�ȗg-;^B�����2z#�c�j��VQ�Z��{U��e���~>�5}�������mBnX,q4�ч��o�mA=�����^&�|uh̒1%O��`�RazS��|K�W )��[�@�p�m��Z�i�=!�C��^���;s3�$G�'R�� ��B��"�־�f)���a�N��BNEl�H7��O՝�~�BzT�BF�	�P>UZ�}��hǤ��b�|�e��X��? �8�P@���XR�Ik����俘��>�]$t^ڋ�%���&��4P��ꄧ#K���ɧ���u���>�05����%��D��2&ygy�C�V��&�����$~��eo4���L@��h_����'�FW��AGC�R`�g���?j���<V���}��L\��a���Gcs�S �q�	�k<K<&`��~����v�5~��N�x.á��9���-Y�)���rf�^�ד�d�p�.��ti���7B�B�܏��	ݤ;��K��e���:"�L;�ٟI���	�}A�����Hzy��˩�,���qm�6������`�EqM:ǅ�~Z�#�����J#3u��%��)��`!���-|+6J,"����r��k��MR��qa�I^���[p:���\��@!�g��_�Q8�ɐk�4��w]���� �wWExb21�0�����S��Ԣ��;��#�|n�Lm�Y)큂���:ؓtǜC�:ZM*�H5�.ɱE����L�I��{?\�j�?}��=z������!�å4a���t���l��>�+TX����0���I�r�n2 ���6_�%�ѥ.��L&oYmՎw����s����[���MƘ�ǳIS��6�D�1scs�6.:�3���"z�|�t�c|�h�Մ_*7Sg!W����4̑&���4�޼������V��V���i	���" �eQ����ׅx�օ�no2�TV����g��]_��ͼ��H41��6c�����>���.�����/�}�_q��X�`T��拏N�~�[q��3�HD�PI��t�L{�$iKh��(�݁��hzcs:aƞT!�\#�f��|���og�z�ݵt ���H�AB~�W�޹{���P��>z�����@��&���ɇeg�.�U��������at?��r��|�� �*�/��G���c���]G�[li��IA~���#�ڕ}�&7�0/�ݕ+x�J�㬍X���c��㋲!o��xDBy��$�(�j&X??92XSn��i]�Z>-*����;�45㐜%���ji\u��
*��pE';���e�ɍ�|`9:'g}Lwo����-�"���@9�,��2J�#�{�QsO�����X�j��1$+��1�Td��GՋ��H����Jhv��.�8214����
ݐQ�w�xs}=�R���E��~��ŗ���� ��fd��<@�cP���PBX�� �ߐ��"x��zb2�=��#�K�m�ڏxgi�ٔYw�<i��J�<E�򂴇z������l��O�����=ߛR���g�����`d���F���#�DV 
�&t�rm6>�V]���])������C_��Z�g�D3gu��2nT�N<.-�s���=�AV$.�E[X�ʚ.(�՘K=�Q���gR*ifCΧL,�~�ÔT���Wf%���j�y����ڳ�x�\<�Z�k"�A��݁�.D����R|��j�(��W�,�ǺU
�$*��)�.]�OL��,� K�$�m�3ba0�]�q�)_�(U+.Y�s,Z��d�����%���� C���וS�	038T�	w4��oֵYk��֋�N���9[S
B�����M]Ͽ2��.���~���'�(������͊���)�?�9�{�kGO�q��5`g�V��X���c&lƗ�f?��V�J)@Z�K����ם���3�xc9�X�FŠ��I��QPLʾ���f��(%�l��f�5(2�P��K�|9���m�Q��NQ����v��	�N��$���sM5~D���vΡ��5$n�]$.M��8p��JÕ֞E�ʜ�a��I�(d\'ŕ w%D���z�nl����Rv�fL��s�<�&p�� 6�T���V%�Ʋ��sN&�4�['
��4� �>�P��SM�8`3/�C�~6���	�'�\�6b���>($m)�f��9�z2)@c�!,�}o5c���
�h�lY��CgDQ��ڦ���I���t�&��Ouz�=��������j�lz�y�i�U��J�3�ک���tR�����M/w��g"�9��T����ж��P�$ɰl �GN�����T�&���}����'���6�spn)��X*,���/�{�Dćri�z�NN%˄ �^#�v i���Ƒ�s ��)Na���c�T;���x�C�%	x��TN��L�dq��\��~0o�`:	ljPvN�L�@I2؏><���k� ��Xz�q1,|?��ӓ�A�R��'ch�*�OZl�j�>�	��gm���Q}�҅���i'@wR��B[m�s�s%�x	F���w�뀳4����ӱm�U��y&�@�B#��nB�duqg��4=��`�y�X��&�B\K�1	�׮W8�I�!���D�e�]KJ?GN/��>�r��w��6��4t�`��
W��Pu�w�i`=���ke��7s��2�а�CB��3��{��NJ]?s�(����<i[��5t��⠴�Ry�Fـ�I���U��H��ї J�kp@��͡&t7c����)�����ϸ�D�P���ǹ{ݝ��/takMw���\ʒ��N�7~{b
~I ge[���d��	�[��7���z
�_�$_hݹ��
�����b��j�f B�^�,M��~8���:���S������; �(z2�TW���W{�'z�(Akrˇ���p���8�~B��q�<���K�������?�dV+R�|u��L�vsk�����6�h�<��h&��a�v�"�ݧ������|��|���O�y��u	��U4u�X�2 !vJ�a��-r�� ���Bű�}ՕC�ƣa�������7m����f�gEu��7-����֊+<k��\��ំC�>���T
̹B��ݾI4�F���ߕ�P&��>6Q���N[�R�+�]�Ii�k��e�ϭb��hճ����ӝ����K`����h�1KS�`ql�T$�$�Y� E;\*���� Rq'� �1:7�O&�o�Ho����t�"+d@�[ #�Ҵ�ﹰdz�^���Dc�{�����Al���aਫp���Wc#�����V�A+0.���ނiG�r[�T�@��z�7��h*�.&WKI���݀�?O	����8�ӂn؍����<��9h��`!���ʬÒ�d'��u���=  ;�g����=(6
d�6Ɋ
�Ϝptv0��E*�K�� G�2�*:�▶�)����2=_Ԑ�/y��͒q��������\A��}�"��z��38�	}��}�Vp�Nҹ�-vn�RqE�����R!��p4�g�#e�tM�yC��Ћ��5���F�
�'�Y��R5���+�	ؼ����팮�g�龕������?]+�/b���8��,�$V����Z8�i�*�Չ5�nc��:�x���C��w�at���i엦�^����
]�<<��4S�`I�_G~ޚ.��1�w�?�W!� �=���B��A+�Z�}�ض���0�sr�2��{�?�v,�0��(ap����G�"g��R��l��b⛳.��jC&�E�*x!��?Ozy��Do����+5���VC��-��e����Q;��f`S%'ČW�+�2:���V��щu��Y�U�+ħ;�j����$DQ gT�3|kDSs}�J塤����D���Luv?�S��_�m�z�����Ⱥ�af?�h8�c��0���@	f������4�Q�4*mH6I��٫��N�(��z�����Ɵ��@���<��?*�@F��`!��^�+��fZRRO�(��$j)DeM���]�p,#}�i�$��8��+���4��3C���8�n���Z��u[�t�b`ӣ,�S3��5����ze�\/-��s&yB�-9�����?�
��2(�a9��"���5X��E�p��l-2��;�n��md�4��S(�}pğ��b�T� ;{�\�"q��|���q�`#��'����\�lX����M����Յ0��O�A5]C˻���	{�Nz��Jw�v�^�K�n��C��9ƒʳ	�1��Z��5O��������[�>�U�Ϳi�6j�#��/\��F,$I�� ���ǉ-�Ŀs7������r�"m��De�c��	@;��p�m�՛KԲzϕ��o�N�Kē�*cM�z��CnV��̾���?4���ȝ��Z�ߩKc�u�����o�c[��ȊB�0{PR�"W�()
r��Ӯ���$߇?D�{��K7<(%�`�ǵ ���[�5`D�LGU{H�7
�2K�Z粫��Xþ���[N�V&B-`�B�2'%T��>�yf!GE�[E7O&U](�Ƅ�s�h��H�8O%�3A�ڒΑ���Hfwd������D(���� X��&J�oRm-�f|�=|���U=*�;3�%�)WB�U�������f2�%��Rt��y��`�<`1�͡���@b��}���I!p`�A����\�0`�M���O��Iӛ�MמTV��F~Yv,h%У�4o�?N���r��3��\�3)d7����?^�c�����^�_�2sՌ�����Yt����p�9�gr�x�?^�y!���ezjZ,�ʷo��tD�Ւ���<����r�d(��ꨅb.%�	�-��?���.��|x�����dH������G����KՓt�m�>����=e��CU9@�Z�( ްN�s�C�R/)���主/М������۝܍��hc�X�W�552s���C�������5�^��R�4�}oFGg���m��1�H��G�����l*�xo�V�}j� ew����i@��}S�!OTY�����ʅz��+�J�������q,b���Ӧ�n[4�tׯ�|{~��< Jt�~��t��A��l�l;'�Ϋ���n͹2J�$j-
��ֱSBe�j���Ch_��G�/�4Y� }�pS�aC��LxSې^�l�b��UB���
���k!>"sHB����SO�*(�s��,�V;�ݳh/�ʉ''�%_i���r�`ˠ渆.����OIYW�]}�@��@dh�{�#��e6�Td[�j;t-��/�<3w��ᒂYwYLr������ 9���H�S�u�̂��q�MV"ö�Lfpq�xO�߅��,Q��@��x�=5�+#_R%)\�O�~W�ρ�6��� �տ��ܷ�u������j�#�KW�p	��S�#i�"R��7���\�Z�!K8T���3H��T��N�J�^�؄��B��7�G|!�v��{�n����Zr�����Sx@�b� hx9�� �`}��jS�B��$�:��r]N�8��Y��� �S��e���ˁ�W]�_l���\�%�Ɛ���w�=o
�с~�4�\2���AQ��$>�Uy�r+#���3V9-�!8�WT���Z��.K	󳎭J�(�=���GL�%��Q�~ÇӯP��.�i�aG��>Y���P��_�xv|�.qZ�& �9̬�+��cMu��K���U�ѐ^H���v�r� k�}�,*m���%�CSbH+��XNH)����q#����-�R��d%��C�·�A��
�k0�s��%k	ң����}m�Q��P�����䏽���pdIݑ��Ј�v{�峉�z�/��>��477t�c/�����H���7�f4�8)����Y�rw��6�����dl��
l�o��D!�����[�J�#RӚ!
�k���-�S�{�<�0B6h��4'����iv�fa�t�82j$��N�5��s�����1Satʁ<���W��7����%�Kp�H3��D�m���C�rA��D{FW�J`�@܂.jèB
;?f�7Gc����;���U�>��km+��+�DS�}	J9�˒��<O��S��Oц�����e�mޚ��]���_�ݠ�����RR���E������E\��
��=}-u��U���	��%p��U�]2X������M���7�ʖ7�A,x2�P/�A�n���u����l�j3���(;A�O��2�k����Up]
�f�";����#�y�(�@)N`���8���@�5?�&k��(�����C�} ���'^ㄦ\����j�i�'s��{��c��t�ɿEB]��L���O��~{ھ�s숏#uw2��g�EC,�������Iڒ$�YW�H̗�W�6�f���N��5 �?G���be���;Ŭ�xk�RLF��~��lΝ~�>����G#YOM������[���͵|�ݨV,�4�V�|w�p;�����}��f	Rw[ܭ�a�A�v�j���J�H�% ��w_�Ez�gGQ�2B���P��z5��*��d�����)�Og�قq�\'�vGFe�'@Tƚ�d���i��X�ӆVU���HB�&��]�e���DS�!I�]��8s��%
^��� ���Q�G(�[dA�<��5!���Gz.Z��ҋpe���JA������,uO��{N�y��֍/s/�����Z��#pz�6�������n(��*B�����J�2M`��}�5�"�F�c�u'3�s����Gx�Nj|G��ث2�N|�K���� U����S!�X	bj��>�˸�m�l{�
����۵ s�\[�m`~���g�Ɏ��b}ж����=#U��jZ/��e�k��k�»ˠ�e/t8�Q��,:]�]6�vQ��;W� ^�L�#I��h�H���u}���_��w��0>�n�R�uSz�������8�R����a��Pb�B�y�;Ѭ�}�7��6���tPbA]{oc��D�R��$�7�GyP��x���ߡZ���T��/��k��&3H��<ڣ0w�q�'R9�
N���W;M�t9QsK-�Ӟ��0y���e�5H�QG	��M�^)l�)7�b��l!M��A�$!j-�D"��� �������Wt7����k1�����F9P�<������1�5h�,��-*�B�
�F\ە�>�L���ku�+�n/A7W��U%���q��u|�$��N@�gʴ��\i��S���x����T�I�R��|hh����.��V��&�c�+Q7�r{Izs�A��9ʲ�9P�So3c.��-��A�R 	��h������.p|?I�y���O�Kq������t2ެ��������m$�a�RZ�\�l��ߎ�\�_���N�D�8����F�۽��J�`Q+�lŽ�);G�>ԝ���z�_:j����?�+����$�(���Ͱ�@�� 7/Hj�}�h�G��uЏ1�˵ �.=Τ��wZ-M�����^�	�(ت൚R�-Ό�����mt�0D]�5W[�&U0%�R�	���QP�w��(�7��΅�����;UDpbY�	�Q�=O��;�"��t��~b���͍�|�HY6{�z۬0
K���P�+�k���tGU���c=S������F53��	e�lq��>m�LM��>��>��wu�Be��� ٛ����8�>��
�gq����0�A�޹~4!�N�|�	I�X*�<���i��n��ts��t"��	񕓃y��A�>�Q=b�1�0N��l�>�q��	��� �CE=�E�j�73m��!��ya�]SR�7d|Ze�`/�W����� w���CӢ�%�"r�C�ꜗ�7y�ʙ�]�H]&�nۅ���Ϟ�)ǋ�.���
T�;�@��e g������2�	�Z�I3z�5ޫ=f68�n#o�ԱX�W�_i��A-4��&MbL2H�=j��w�bX��Z�������=��!�]�ǂ�[˽��Iޗk'̄�y�/�[�b�7z��S�+��(g��W�/7�n&�Ʌ���
ME�k�p�)V���r���� w�G?�z0E�a�w#�����H5�2�#!��t[�2�z��ܔ�<`A~E ��O�QM�[�c�Q��؀h:[�B^t:���ޡ�c�]CA5,����q*W�
�ǰF��h��{�Ak1����5����l	�8��ճ�#]��&!h�H��;��e���QƤ�ݤ��e}���.x͓u<��A%j�#���vs,엾Ҥ�j������mi��eg�kH���X��7VaAL8"��NN�� rOBl�;3��b�f�&�p6�W�����7���Ԑ��23����6�a�v[�Oy�T�#r�2�U��V�@��𞪃/r���e�+Z�"H&!dѓ&�Q�;�m%�ޮ��� �3�k*����e�M�a,��Sw/V���,�1���6 ��K�d���7�m4�{�L�l@w��:}��������\ď@�mz�<rL�U����Ƃ���o9�!�b�<�K���E���T�����hBNR�Qh���ct}z���ݠ�h0\}%H��@)Uz2����q]M�e���6��0�"ՠ��ڃx���3�-j�頣Ȩ؜�_'K���O�锅�9j����C]޴,~"zBs<qᢅ�,�]A%'mNm�1��Ԫ���԰x$��k�4��r�f�zH�����	�L���������Dq�|�S��C�i�DiE<����_ҥ�z�!1C}���dj�,x�zu��a�E�����KC���M�i�/dJ2H�j�u�h�M7Xv����k�]�'�L������i�T����INt}Ba�p^i�0
n"��Tu���q��n�y�7�П�|RK�+H���O��O͊WI���u�MX'�V�NB�ዺ��j�� [�
�U� ���{"��Jjy�|�Mc�!&@�*�*)�6u�L3R#/PY%���Q���S&�(n��veLx���ʡ�c��t����d8w�ļ�Mਾ�M�s�i�.ݽ���mMǐ$��">���IVS1�_~5�>9�;0��f8�@�Ee��|g����??
��'�Й���0�vM1�ȔC�a�?� [��c�Ua	~.�f���Y^��b��A�	]|�	�/�olj�z�mj��~�!�Ѭ�Q�LU(;�'i���$E |�Q��>TƂ���MҚL����n�u�����>���
�h"/��R���po�؜X�=�ב�"���^M �C�}�o�7�`����:t���	����ep�e4�OzF�f��䝐LL���|r�R �p��i_|W��Z�xh�\D���5�t4�M�W�n�ψ����R)3��"		��giZnѽ8{�&�+A��l�K��='�|\��s��o���ҕ�-!�B�u`�gQ�o�x�R;���࢙��J�Q}���ȻH����z%���T�S�������B��#b
�ݺX{X�Y��RF�����-]��P��vã��*Y�Ol��f�0P�t��؉[B���Z-5�2�#�
J����[�!I�o��*�[S�ݺ��5.\�`H��b/\�	��`��^G���odw���F~g͔)��'��-�����"��c�C�8�^���m�;�v(�W��qw��v�r}�(\w�1Ջ[�qۼ+��%��o.��%�.��
���I�y���R�aZF���ۖ_�W�-��h6o��|s�>"�v��AT`�,9

��).���J�?)1F��!Y�y:���Ӥ듒�9�ȓ�/#�;6�Ȏ+DW�w���e;ଁ(�q!d8o�1i���y��%\�/��-U���*�?�UU���\%$HT��3�P���p}���J�|[
�ql���|�[� �>��y�`����0@ܡ[F������p_,<u45�a�L���>N�)�"�L2�Tʏ�!�^��}O��g܋k1Pg����A�հ�W�j��z����t�/����hk��_��2 ����+�-�pE�`0�M�/�ۆF.��N�G���+�M(v�W�.�����o�n�i�ʓ���k��`��י���D���Z;, �d�'8��r��0H�R��M7�o�he{��L�8Ĭ�Z�^��� ��d�f����>�(0&��������,�⛆G�mor�PEAAh����X� %u25t��(��%�1�(�E-K�d��(j�ll��Xɀ`ysg?MI�w86l�g�w��|'�Aau�����U�7c>)o+�ʞ^���)޵[Wcd���C?C��)/��$��[%�~�G���J�ZH<�˙��wk�:a��a}.+��%/��o	��N�BI�㼇>lCQv��t�I��Ɋb��	�R]/��y���$xA;����G&_�<�D�S�ˋ�"˫,ˇ<����t�i%�2���w��'&���Ò�	&�h�&c�NQ�0b^,\϶O�c�^�XhJXZ�>z�bOOH6�B}�@�A"�h�:�$�7����yq����b�x"E���ԧ��!{F��P���C��*��#��k�iƒT:Pz����G����g�!�!S��ဲ�*/�;�Ύ�JA1C��w�x����1̀� 3��w�J��ܾ�a�R�OS�1w��=
Bpj-��������	A�Ec�(�-Z��Q QQ���P��I�4
��p#���ǥo�ۃ8l��V���U��GD��%*��p	�����A�2�*�Z��٩�`�_	.g���� q�V������ �6��CԞ�zn+��@��Od�H��Y��ˉ�G�:�(���)�C:ғ�D@7����UU�����`zF�J�W��w���bc0+���`!��};&�NB�J8��ȜL�`��n�23F�V����U����{2���2�Q�]��iD�]��=�h��W?NkQ=� �Z����ێ��ח�H����A�t���X��[P#	��c�j��jA�O��u�qD��x�� s?�@��-s��T����ȈO�d���J����ف��yE���(�� �1z��@#�{?F�oj���@b��8�v�aV:h^ae~�o��֯�ɷ?0vh�1mc��飀ŀ�=�d"�A�;�Ay'�iB�h�/�Z��(���G�r�6��BR�]�ʆ��Z`ovR�zV�M�bU燆��M��d��n&��*�Ƈϟ��ޓ����O�߬2S�uy=u�b�)���m�"�T�O��S�C��Tr�q�F��`�qt?��~����Z�E%�����f�5ϪM�w@�/�q[�["�}�[��Ĭ���l9L��󹔘0�d����g8hf
�����~�L�\X�K�
�ql��"�ťSp������o��*�}P5r%\�'��I�À@�נ"b�$�������=ۻ������sf0q0t�V!�S��M�'��x�F�K��u�\қ�>%؉� �&|<&�\&%g�tA%��T�:��v��.7pN�qyy��R`�k�f!�
�S�s 3R��q��z��l�bC��3 �O�CV;���'k"rO�h�E�W@R������T"'�!?�0`_�=�<���{����y���K};�Q0�^ZE�D#\�zsqtSg;�$�R�5�Ǣ;�6�x.<#��ѩ� ��LH���s6�J�eEW~��ȉ��'\�+^s�To��.2�?9�v'#=%S�ٞ�E��w��(��y���K�R�ivh��[k�iˋe����s��S�ڥhY��x�f���aQ�ZNb�/���F`�kr���yr4<�:Ţ)ľ�����f��Kh���=G8�Yv��%�V������SY�μ}��fz
¨:F��\4��>��9y^y�HGO'�%2�cS��0�Aһ��9�%���W�">�Ť�ᩃ�2 ��1�d5lZ:
��^���i�
bX[���Pc%0����l)�6�2���,P�FFD����RX�>���c���{�
g4�U��F6h��`��ե3��7Z�y
ڪS:{�y���r�ђn����
O9�͋tg|���kx�X����3���]��K�����7�ho���=x�v&�ɒb�v���;u�rQ�9���Ț�)��*��MP�e�cg!�5,����/�K�~C�{�����zKp�x	B\ф��3� ��
�^�t�j��� ��N���}
�ֿ#G��{�:GsU��
>�!�/�F!��̞�7��B��3j5�Y�_����Q�FiC���B��1������%�E�ՠy�{���������N�ok�ώ[
���!�b2Yf�N�wz�[i�7�:��ޔ�Ȟp�g����O��j/�c���H������t���Y\<n� q#//L(h�I��&��L{���C���N(��Wp��f"BӰ�-럑��Ϥ!m��D>��Q�f�4E2 ��.׻Y��K��#x��n7؉����C���d�%����/t����V�ר*��H�TiK�Y�|Lˣ�@�X��8$ +�9�yа�4+�7��֟�.�3K׌�Z%.oLg�}Ά{�-�� Řs��l�dE��|#�	R�I����]� U��cϊ,������؞Έ)��@�f&�IWo.��������ݨ�j�/�(���}!
��7�b�ȭ�ǞJՉ^���σ����z��>��O�3��4��	���	}bs��q�5k%c����f����v<;��(���0i.�"���J���D0`�����9�f�-(n�wD��=�񐚥��>�Gc�f��7��@�t�#�0�7���[�R
�|9�`B�{s����pB �-�"�v�SAt|vg�1����� ��s­�[���ܹ��4�h�S��/[2�%u�ڪ��R2R1x�O�b���A��h�ע]*]_���`�cF��tF��k��@Ū�����s�,@�F�uo�už��3�$�EN����Go�#s�d�O8�0/�����-�&I��!�$cM��I۩x@kv�b[�/������*K_Co����ķ��Cf��}}8ˏ��j� �n�{��e��$M��9\d�1�{&��ry��5
�U9+�i�u5�(�X;k�Ԥ5TAqj��b
{e�ܡ�9j��s��{v~P��a��V47� �;O��3����k}���5�rNc㐦��p�^!��S�ڑ˦���,�&���Z�$���<�S$�ށS�{��:,<�$���A�TE����ޟ)Ej#F�)���G>�N�g��^L���kC��@|ѝj7�b1�o���6:~cS�����A��(3@�i/�`���Ȃ�����p�PMZ�6~8��J;��0Y���o7@ɝ�LF����G�4"�y�0�^~0��­/�����냭2��ݻ n�U ,�-=+f0Xr.� X�)�$�}�ՠ@T='��+מ�_��$�7K��gG�6v��2l@�r����XT����ҒΆ@5̩�����C���Z��n�Jæߤ4�2r���������֖dƪ�/WJ1Je�~{�_��S�4/�A���1�sg�G���a�3J�<�X�|v��k�����./�ZQޏ%��EY�`���3�֛����v̵WwD ����}��>�q}��-�Ë�+!��zJ����S|�v y����ߡ��9 s���4�oZK�
�m�Y��7O�!"�"@���
bW8vo6S*�E�����Ъ��m�N�ٓO[��B�Q2��a]m�r��ج��t0��0L�"��>�{g����I@���D08��9o�s���s_x$%�����&V�������UZ.7����oL�j�X_��I��^w�v�|2d�ɛKGRc��Ͷ i�����,҂a�nd#�tU�4y��˩Ѕ�P�h����0�>�\=����t�\��YF���.���=-^� ���iN��?��*&]i���;�c��Z�:��׍��)*�oD���B}G����� V/�d���D��`�@��Br�ſ. �c���?�=*;C�C�d9B�cu���<�~��/>�i(��|�(u?J��F&��I*��L�����Rh���3���f�����`Q2����/`PA��k5X��*�D���K��iE%�Y	Ä��>�ak|
*]�$��d��Kc����q�V���;T}�.bµҏ�ړ�b�9�%c9��#8WM\�pE���[�
�6��J����*T��\�i#�`[ԑ���<&����br�O� �1���Q�IDS�ύ�y��e�<G�ɟ�0�Ѥ�Ϣ��T�Pjq��z��v�~�x<���5_-�o �El`���U��PjT`O�%Ϭ7,`!�x�Os��]�ן�(p�}��RO�p�ID�Z�Qt�Z��fAހ�n�]?g�t�j���/�=�Z��
���ܴK�`�5g5��;�X�`ЃT�=�@9$a�f���H��l,��X h�h�����+'ȹ�Χ-C]��7V�*t�4����W���'×�I��3����i���R�J�-ݭ��/`/�Y#چ�����? �.�AnKQ�@�"�~�D������*lzҎ��~�����M��?����t��Y���.xO���@�IŹ�]C�M���_EL8��D���N�F�ON\ R<�'Sp'�u�b��<��0�,'8�*R���ot�7�	�����eDF����R���y�>���gJ2���m�'�~���u���Z����E߿2E�z���1�b�YҰ/��(`���P�#�%=�5� [�|�	��?>�S�/3	�j׉|,��-�5eW�T^��7�9t�qο��t�z��D�^��&�(�y���+=n#�q�Ig~n��7t��9p�OK��9G%[h���6t�O'�{�)r�������)��*S�D���ݎT�of�<�X�Y��G�\�#z6�:��+6n�n8����׌h��7#��7�C�\��P#�ny؋�'��[pj}`�#y(ǯ)�*{b�d4�sgQ+��n�胤�;���}��1��տ��O-��<�10���|̭w1����Y�@�ֿ��.�.,�:GV�O��z�	v�'slp�jN*�qc�:ܟ?�gZf>�]�@�s�*�f�1�J�G�~;��y��h{�ٚ�}�����Ǻ)�b���-��r��p<��Ε��ۡ�l��2�Z����n����n[��%�\Y�>T�.�'*�Ra���hm=5x��˰K�o�]Y�o�)�3{}D�`��!�f?X�1)�����'{@=���[�Ƞ؀�>=-@l7v���[�_b�G��]�Zlf�nk��2�����h���+j�h�����n���B��+鏺Q_дS����� �O�\�R_@�񺇬5�������bs)�iU�sR��h�f��de����c!�����6F����}0nY�z
Ǚe�MW�{��k��Q��b%�� m�����yX׏�BI�o�y��� �L�Ld?S����؛���u�t��qθ��eO�Ad�N��g�1С/�+�%5��f�GG����gƁ	��/���\�=�����(�6���ذ��i����E��%-��)}d�)��8fIU�FE�y�&'���D5걦$5U�� �{�z�H�O�iOv|�8�%��+ߦ�{g CD�Rt��rK��<u/C���a2��,���;��n�(b��gh�P��׊M�)h�H���r�A���%��뚉��]�@�]��?�) !��y�W��r��p[y~6��r��em%*�1B̐�Ɔ�x��]���q��uy���rhܳo2L<����mQY��4S�K#.����<�k����O�����u�t�'�
n䍋����7梙T�x����Q�'LtM��l�ܮ�#Z��;�E��G��^�ڕ+��}�+h�t�lE�D�n�h�x�(�>:���(���G�RL��|�t,$]d�A��d���k*j��b�O7K�
Z/zg;��f��`�x]�,���?B˾���m�R��i�~Zyr�m�~�|�[	��J��|�*I~Ӱ���������g�mS})���O��@f�?����1+�^f#� �q=���11�~��:�;���ZHXw��[~���b��{o)������,�ar1�lp^^D���CB��e��x��cz�\��M� yƑ���يJ{X[O/����W_�5#݅�����9Z{:?e�����I]�j��)V;L�^d=Ac�s\�
UD�my�����e^!��'��Ϊ�패zXV����.� M������XFo��Xj����� �PPH�(�tL�F�iF�b���Q��Q=f�Mr{h�f�K���d� 8�t�9ȡ�r��3�Ն{���UG�!az"��.��C2A:�g�+��웭WVc��G�q����5۱��
�ޅ��������1�����иk�����!p�!����8������;��tdD��1lNtPCP�֐m�5q]����H��Wԏ]�9�+^w�&�z�\\gz��!k�ReXZb�w�G˄0XH�[�����4� &�V��>��S?��C���U�� jjڏI�8Er��AfG�\���j~�K��a˔���E��H��]���qr�T�s;LP���}:C�j������hgz�C:���k'e�UCM����,�Fj����\˅��2�ڮ��(_�)��"4�
kZ��� ����H��@�w}���Ӯ�%�2r]�h|a��(ΰH�>���������>���@ʝ�mѢ��(p�o��vˑ�ɟ7}_���cX��_x/AS(['��L�_����j���eJ `yW��L����Jc#[����O�I��2<���(�k�3r���ӳqL�M���	\���Ӟ�V�(��Se�pY5=�7c*٥OZ�S���eP���G�A�H{ˁ�4�[9��<p��b�R�^L�0��s��NΞ���;��S��"�/b�oSC|�q2�70�(ݥˎj��Q��[?MYCY!9�a2��[c�l�1l�1<��+.��kK^+�,�m�K���ރH�.��W�^<�����2I%�àI���{�=��;�t����3Q�� ��6���7�V���]����f �!zN~���L���Dޭ�Gj~]��Q��B�=p��Ө,ߧ�SOZ��ؓd�� ���=Az�� ��P��R�H5��G�6�7Uƅ�jU��=Ԝ0�>�����?�E�ag�̤e�>�}@�p�㼱��ݚ~8��E�`x�p�����q��r�E��K�kփ�f+���s�����v]�1�)q�cO���e�
W�_��ށBf�u5��$��u�&�0H8��Vk�9��e��^yF+#�@�aR���4�(� ��]T�X�w�� 1�����B�
y+�ˎ�M���� �\ZcGo�[�M�))u��j�<��l����2m��U�����dp��z4D�MR	�L��X؞�j���~����v�0A=$��lA��!��P΁O� q	�����-(j���	����ʉ�s��,>9rF?��7���I�`=��ٹ�FRgf{r�ė,��<mq�ō�Dĝ��,�N�~�O��=^���Z�Y,a���FD�5 p�����o������r����	����2��t$���E��-���/Ҥ��)�9�+ >�Z���}��3���*�ʈ�I;Z�6�<7�݁��G�ҥ�`b�E������Ee��V���8ꎻ�퟇m�uD�������M����YT��|F~#e��&�k��9��tF$e��0��$Sr�΋��t��f��ҵ�Ӥ���/c38]X]����Ki"��A�����tN�z�ݯ�v������fs��A5nJ�k�o��<��B�:�Ԍ>	C����JR~� 8S>Âe�B�#������l9:�fUޯ'̖�B�/���"����8��m���_���X.N������O�>�\�����x~�hĴ����9�.Y�� �9:
%�2��/�)��(gt������x&)�uL}%��J�ڑ���("n	4>zY5q�^�PdWK�q��ޭ�M$�2>xo��s�@��N��e
��� /.ܖ*$�$t@����y�������37�|׈[�����,�MX����QN��<���m�b-�)������6V������LE�7�v�L�thI{��������Q]�6g��V6˝�\�m��,��T���n��������qَ�xJ��jVӘD�^Pm�QɰZ��)֡B�ݰ�X���{~z�����Ü�	��������`#jNY���6
f���j�at�s�o}��Z�q^����5�z�؅��#]��vļcdŢ��df���O[����B��HFN�ߔ5h�LO����餘�?��U~�����p->�كH���4�#� 8�Myqd����Jn���7��h^�MH�<b+bWm��C�2�gK&�� ͂��FÒ0���~	��*�?�����w+�ZX쥈�xkTG��C�J'5��:"
�_=Ox-t��S��*}�Y�W���9�ZP���p��� A�[�v_�d�2W�@�4!9S�r��)\�ܩ@�z8H�>ϫ��W�:�E��3���z�����R
��`��B�M��#�$yJE��}/{�7�U���F��Pks=gDd��'Q���Sta�'�r|_K�I&qq�_���o���uI���W� c�ˍ\Y6?F�̮�;�-�Y�~1P�1���߀���=��A������9�i\�����m�(���E��W=X ���v8
_�	��T�W�ٕ��Ȍr/�Έ�D�1N�q�^��p��6&�� 	S'����rV4>����Y�����jR���GN����+f8�u3� ئ |#�dn��<?���w$�I�J3��@�ċ�2V2�(�'�����t6E3�����6�Qc�����鲘_J�S�Iл�l��߲���^C@�?tڽ��)ϒ���Lj�^3��o�f����7��P���5/�v�9�p@z��ǵ������6Ѕ�$$�0;��L*�֑h�D�G����<�l�<@{��x3J�x�jgC�J�T3���l Y��ck�� ���<�������q�aqR_�MjJ$�L�$�h��X�6c��nMӶ8:!KՖ&�0Q���"�ӊr�/#8��vo��X<{ݼ�6Rd�i�!��Kǋ���_IP�g%�'�]�"���"�Qki�ȭ��ؗb�>��A���4T�D#*U�K�+Ө2�$��g���W�����o�u4�0s�\�~O���������l��ʏ^&�/��9E@��EI&޽�GS.J9{��~s�����(�r+�
Cd���Q�e .�;?K �3�#E��lEnh6�x�snW�yBw;V³�"�#��������r��Ī(�N,�Ι�'��a�=Z/���պ+�#=�`OjO&d����D��^����8S�>��Mz?��r�>��Ŷ��Z4Q;�3�������{��S,�]	�Y���n]�z�[�_�7�?�\s��٣j6B'u�I �I���(0vVPS���K���Bps47\."��C�(̋�/��Sp�v̤p>���Un��=]U<|��z�����?�A*��2�����R�T����J�xcX��&b���(�n[k���6�?�4SF�jH�m��(���t��+��O��7T&��k��Z͠�J�u�m��y�����E�1��M ��P]�(H}u	F� ��E����L^�O�h?|�d܈i�F+�U���+nV���0�1�~��������G�|O��t��7z��]u���s��-ȇN��Br���g�f.��t=�u=��Ys'��w�[�E�/��J�kP�%� 6�D�/xagGg�R��{����(�y}��)��n���.5.NV�b�s���,�פ�x���Y)�W"�������݊�ݞ��8^����/Myӄ
�¹Y�J���guƠ`���X�e��2��A��A(��,����֗�HԞ������B��5���[f��$@�V��A��@Y4�pn��4� 7q>��䙧��k�	FÏ�8_�"��?�0�#.E8�\�<�&u8F��u�����`Jb����`��/�P6��d�J����U&�8F9����m�����l�e�l�P�n��R�l&����T�	6��$�*���C˓>q� Q��9�\C���� �&M����?bcj�H�ԍH��v|G��x>���m��Zf�Z p�$�RN�V�W�%w!<l�ԑ���[z~�m�djan�����m�C����/W��s�wm��L	!��v�UKyc��)�Be�Wt�Rk����&�O��Eyx#b�d/�'��4~�=�[!�+���Ʋ��a}͐��q?ᢝ�0p��.D�:òO�;������>����Do��L&;6Z�P�qp�Is$��@`06xlA��^g5���ٵ�����+=� ��0�9d夷��u���55�rǎ(�6������S\�IBiN_0�ĬIf�n�d�]�v��e�dB���Kڋ��'��J8����D3��(�-�	ʪ��&EXy����#�ʪ�������ᗟ�_��.�� �A)-�n
�~��������:"[wӎ��Һ�)Ķo�ˁ	�$~�_~N���+���}�=�yS�r�*�Q3���|��%�s����ӵ0��-��U��$'��5��þǠf_�wh�ˏk0o'г����;K{�HM���k���⺛cc(if#yw���)�&o�{=�HF�7���Cx(���px�=��3�
@Og�-����xd����}���ڛR��i^g~�tT��YテȮ�A5����)ƒW�pe��k��j��o̫.B&$�e_Ɯz�>B=�p���{l�gg�O�
4-�v0�*��Oh3ͳÖXO��卙�s������ %]�tH%-����_�n%�*¹o��J��eN��\T���z�C��Ņ�����B����ʩ�c�𒂓F�V|Ѹ�s��хꌆe���:�Ug��V���h_�ˣ|%R�x�ahⓕ.��W���[t	�ۥi�w���R��ڹ�`�:y<�GM�_p\iQ��N�dEx+����a��v?� g>磻Q9�a�����o�p2C��!�J��5����V��o-�S(��p��	���8g�uBJ��
�,~ӆ�_~�Y+]\ �]��_ڬ���1t���\ ��a��b�~Cԯ�hl�T������ċ�޵P.��k�gp������R�HQ�+���	��.��T_�D5Dc2���&�����\�-k�ENԣ��/ �K��H�vs�4V���L��Z=�������"Q��ZϮC��~0i������z�l�F�,�$��3����
�TȺK���2���W}����M5�	ˡ���V� f��Kr��&&��8@�n~���ޚ��\S	F�k�TK�[�oEz\��� B=,!��dA��:O���pCz�'s�*�x�x���r��(>)M��
��Q��E�UT��1x�yn��'��uY� m�M�t��q'ts�]lf<��l2�xKlÛ\���h���"H���$�,q�,H�>:����Wv��y��� tUec���[V�1E�Jhԫ=�8�Ă݄�
"�[�Y��8OT:1����!m�/��I.c9�\�C���hiCR��8L8����4�;�� �q3�V'XWC	Nu�8G�0{�.���Aҏg�h �hU�"k]�����6�b>G������MAA$s�K�x��yJ�j��Ż��4�&>�����U�S�
������r��b����ua5��<P�ȭk,H��Lr�ܖ�����ճ�����8��ϓ?U\��0D��A}��ñ�3�F���lՇ�Ȕ���X�L�>�#��Κ�XJ��D��.M���t �1��3R$�t������7:rǓw�)!A��W��U?�����	?���۽�cgpJD����~�-��4a�]V���#���/�y`x�T�"8Bg}*�4N��ܨX�y%
����������.^���9@�>���s��&��� *�򞟶�߼��R~�u`�`+�H�z������7gO��$×����ނĹ���uF����=:�bJ1�?�� �L��&H���My�P�:�"O�Wd����6���+�$��"�͂tl\'����	�c���=�%߰y
��	&\��B�m�qFߝ)���t-�S����#8�H���l�����}���x�AN�H�x���g�T�Q7�^���t~y�c���q:+�d%�~�=����NAP{%��I�H:�*3�I} �`�<y`}%:`�zp�#�HR�B����۽�8��:U8��蛂
���D�́,ݒ[8����m<�Y�l��ܳry��f�=nw�0�O.}�e���
�G��+�0^4�����oI��-�ĝ� @|E�n����c��? ���P�ȡN2k�`Ϸl?q����v;�h�r-E��
b����X��ZH�h8�\ ��3#��R���V�cp�_��?��&�+�@�s���a�<�4�t�O��ܧ==�mu��K.��F1H������ ����j���5W�t
�iV�64G��j�XZ>j���
�4�m�$�=��z�}�ؑbV2E^��8�x��y�o��ŊNM1.7�iH���z;���.�pO�H(m.?��z�~-O~�ϯ6�őe��G5n����͢��#^Y�r�����Lmp����+v*��p֞Mnux�)������V�w� ���X�L3&��P�Z�Y���
����ȿ��+06���CA���B���_w���o�V����Қ�v=�슅�-[���F�a��L[H����W�"4�qߝ��G
$͍�E��>�"��������ϰu@�c�2Y�j��պ�bJŃP6��ɜ鰵�	�5Ҵ���T��aW�v�C{BS-�o��!/�wly�E}���3�j���oz�e΀���CD$4(��Z +%lU�fV¸hJr#�ȇ��n��1�dSڛC��^�s�$�¢QЌvj?��}�k	
Ƥ��ŵ�؟��Q�s#��y��e�E�i~z�� L��VA�CB_(�� M8x;i�r����"{q/�֊�Qv��19�Z�z�g��#�]^�T��v��� Q�#t�F)1dڠ0H��kJt�'d�]�G@� �����&��Ӷ�o=q�+t�w�+(��%{$�tx� �����b� �ƼI񡊄�gU��MUku��:E��0N�-b���qmp�"�i���51�;m8�`��m�����T��;�*����~����_R���g�N�k�tMlG	Nzqe��us��e��I���
^ɸze7G-V��n��1y�8�&?'��9��i7h<�J�����U��n�O`D"��e�!�^�̸N��d$y 	�|<�,��
w%�@�T"�r5���P� ���k���[�]/�kOG��@�8�^�Y29����FK��$��d�M�/X���.u!����X���9q�uX�w�	a����D<������7�J~�OB��z*׈��CA�Glj����_#�[+ �p��Փ�Î���+��iؤ�ak�։��T�:e�#�hjG(BV��W1�!�,��hu�L�?����?5j҄"��qM��.�+r�O(��>�p��=��j_����k]8G��Q+���1F�Q���4�]��)�~z�򺀫	�QE2��) �s��4�p���,j��򈮲�9W!��6�5��ؘB)R��8-c�D|B�k�z�qߞ<T^��j��K���`�׆�)>�b>v��_sl��m;��g�fO�>�\ʜ�co�7򓒰K�\	��۪6��!�f���Sh�*��Im�~�T�Y�2�*����ƥ�<X��v��UC"@"�M�Z��"�� b����MS��=Ɗ���`�lٝ��+ 	Q��	�T�M�y�,�A^�e2澫���u��:�y�oPWP����l�x֤$|K���kة4 �����F��k�K�.e3�z��;�;��~dTU��睨Y]Y����|<�T��^/��$�n�,=��J���@��>�W�/{�`rq�*�V�r����.�hv,���^�_\�|�	��OM&�g����읤���
%� z�#f�SM+���-2g�b����g�f)��V��En�EŃlZ�/,9�k݄�o5��&9./M�{O��b��^Y���'�;=/�V�u2�F�Mtmt�V�h�#3���!y�&7���C���A�7JZ,���,4�#*P��^��,�~o��4���eG��vZI�i�l�k_)�S����v�	~1߯�Uz�r�BVaǺ	0j�IJ�%�.��|lf����m�0�Mw�W]bb������x5���5Œ����+��T�3�3�����j��1����e��<�cS���H���)�@�Aܺ�*�D�oݫ��c��	Ws4��6�j��q�3�%�0	�v{#��p����8 �Yh�!��u��<������_8��Z6��e��:�7����ˀ���DH�փ�3�f^2�.6?��Y��5������{g��{�z����K�\���W$�m�q�b<�J��x��;�w��W��?�feڜ���VU+�����R�@�4���7<I��(���!�`1����|=��W�%^
�$���j�sr7�l�\	,���m���!���JmD!Y%mO_�"<ȹ{lknl�"q�2QKVj�nɚ��b��!�
®�!����K��P�k���2B*��5W�R�C�>����Q`�B�G��|��@V�x�ٖrw�{s�v��G���"Q���6Y�|�t�6�w'��z�		�L@�hq7K>���΅���PCKDt|JeNzJ�n��7&V��¢�K�B;ݺ$ ��;9L�����B!A`A)z�������K������w-��s�*H���.�(.�^H���H�_��G�>��cP�>Ҟ�Ǭ�-llדl9�T� ��G�¼����7� �o�0&d�r����g��B�=�W��J(R�9LK��k���s�b_ʡ$(՛Q��M��1-Z�g�H3�`D�.���{���d��XBvx[����
d(��i �e3�iD(�(=?lu9���fJ��0��`<K��Hm�P�+἞�'@Lڰĺ?H�Wtq\�!w�+7\��@	��W��O{��"�ࣕ�jV�"�M�5�ϥ�O�vN/x�Y�b '��$�I�G��v�iCR�,�J01#I��Hs��Lj��N����}l�,Wg�3ǜp�޷m
�Bɻ=���1���)�A,�2�d��Ȭ�B��b��ы��o�6Ed���L����������0���p3���v%����U	�;������?}��k%k�X�3��,�Ў`�ˡ߶g��=�\����⟟Ng��vm̙��>=�톛RN��8��2ct]��S���iҰ,�����]�5��5a�� #�q+՜��x1?d}N��
2N��Dj��E�
��e`ߚ��U�(���8=����H	\�p�lg#��E�����n]tJ�ҭ�gO��5���c~��_�\�j(*���[��dn�r�:�jg�.�Rq�}t\�ώ&-@���`?+��i�>���B��쇑��%w�D���Q�w?��
�JF��S��������a�e�/e���U@^����G�ч��x����P�V��Ô�%=�''�s����ݐQX���1����4M��7�>=�mi����d�崳d�(��e�ri���p����LG(f9Z�!䲶��x��p��jM�J5;�H��%��+z�UK�����ԞDn�rq�.��~�&Ą�E�
�MAx%�+XdjBxc�O�A�h�A�+;��8��o� T�}k_�%J��Yӳ9�<ҵ��4��o@�эB��Z�5�ݸ�*P��eN93�G���*���1�|}���TJ�[&��s���?�X)�y�F�;�#�A�Gt�v�'h]���>㦰K~�^]�I�
���㺒��K�bq��R�AC+�b��sm~j�?�<U{"��>���
$-^mg��sXE���qW�b2��N�s�-R
ܙ|�l��/��y�I��Sb1oiQ)�'���jw�[˗k�'�NX�AV�:�R��T\.�weӀ���-(2-�z��seKI 9�]�c^g�ȱ��S��$�e}Ur1 Oؼ�������Sc�[���d,�(\�������N-�V]D9�k�m^���f��ݻJ�����j��m��X�� 9�@��#�­�0�o�M��6ãbk\ѻ�M���z1Vdi]v1�&�	 ��I�����U�P�������M��S���UHz��oKP�̭�xK��Ϡڠ�*�>�j��XW��"[3� 77��3M�f-��%�%-��'�D�44�~�A��J(-6�>��E��I����;�_��[˦:՜_e����s��[�]:�#�I6����)����%x&N)��9z7V[�aV�0���7lB�h�ؒ�2[�IUЅS��w��b��߆r5�{O������S ?�׽�dD�L��sVk1M(�\�S��1�ͥ� �?W7�#H�?�$k�edY��r�8P��z@>2WIc9d���v�˩Z����iF��z������8�L8{	&�h80w-�MC��In���RS��''.tEG�
Pd�!=;LU��)������o1�����l_��B˭8 ���~&#��.@�惸�~];�n��������
�ս"]�C��z�8�;�����q����$��~���Bk�Պ�~S��fԩ�2�M.�
��WF/������x��$��⥇�%�oDy����b�3��V���{.�AD���j�L'xM�n5Z�'�Rd~�ԋ���e�E�|CrP1R��pE��W���ҏ�����5O~&O�]�5�}��_����c5�"��~�
9dmݳ��jY���j��oxdZ�u\a�)Y^D�Ȋ�e�k�Kf�Fz�p@ā3����p@1�`����@�~���p��D`��4w�㣬D�W�bLG/Q��k` 7�������}0����0��ؽ��%P2	j?���ń����_��zf�{������{Ll�v�W	OG�fj�-��u�8/O�u#�y�]���*��g�C��`�kG-g7_t�Y�~V}��;����8��ˬ�@K-/���0C���t��EhȗF�[�/1&)���lQ)��M��u��~�T���x�1��9�i�"b�я�̆�y� 6��r�Vm��c�g4�#�Ah�A��F���xJ5��4���A5Z�TeUtγ�ȳ�H?�peCt����8>�̩��:�������R5Y�@�H/v�-���]� s�ʵ�C�-��Z�9�V��A0��kU �u�n��E��w���]�0|+/���6��!��=�J^Ń��jUU�:s�GCg�Pff_�7fl�4�Խ������� ���%��2��8}���U�ⅧVS�ۃv1�,����؀�$��诳� nw��k@|�|1���g:�SM�'@*�glxH~��40�/��43��M^�y3C�4a�6Kz�$R�խ[���N�h���T=0mP`\ca��և�؉��g\���G��Z*�1�Čﯴ�a�����N�#�LN��E%n&��l��gL��9��p=/��k!��v���L�͡3��Zz�C���Z4T�����h+$D&�����F<��
���e.j�b1�Õ�uA0;����l!͐t;*����mwvHѓP�b�yA`���N�e��� ���k#��/߫|�qRH�����1�p@�wH_�&��$�mm�);pT[ӄ��~i�VF.�&�XI��K-Z3o3����f9�m��`&๏�4!�f�+T�XP�a`1�T�%�xբ�|�r��<Y8[&�]\�~f�EX�j"��0?5�b�4k�l�� P9�a��7R����z(������&�c�nﻩ{��|Sœt/�qsH���J�q�w!����
�*�9;����Sk1H�;Zt���򜎚��R%��!���-T��?�M�÷�VZ@�|g�sTP�a���4謦���W8��F�C/a��7�v��~�P\p��z4U4��M�1	��ܳ��l�毕�2ȭ>���m�߆�������_�~y~}��!���4�gR�8#��])��C�fγvx��T���u�;�w1I����z�=�<����p6�%� n#�PU3���]֌�� �n��-���$+�翭��!D��'B��y�tS�YG��}|36YB��i�����K��車4#T;o��Cg9��!�a~lY����N��qf�}��;�1U�o�m�&#<�[I��S��y��)K�wrs�LG��%�(H��9��#�M恇�f�wY����/!3��أO5�0k;<"д�����-��6~�3�SٵV�lK&|����C�s��J�g���Sq*@��Yb'\�"q�O�|7�%�E�(i:2��?l���Y��:^��r������s�'�A��~����R�g�ѩ�渘�FZ3�h?��xFG�?���S����-�*�e��٠��ysc���P����t��`~�bq�n�1}�`s�a�k���ݞ�3�1���	*G�p� ��2�G���!B�bX��+�Q��-��	M�J/�
���|?P�xy'�k�����\��m�AZ��!���ӳ4״,���3eF�V�B"}��E|MN'�?�ý�f^�^Ft父9*N�����zd���T��cb���OLrd�S'�ߪX֪Ç�xl� v��B�PI�[G�V�C7��
7����M�������Oh��x�b�V�9%�V�J��5�#�����c�~A/ђ����ƍC6K�7�w!��pvK��p^�ov���p�t��,𷋳�+�Ƀ`��2�z1�����Ԃ�H�W��N���9z�w{��"��#�~J�è�[]_��p��97���fk x&>i�~ �B��j�
�ޕ���+�^���P��]{�<�\(�T)�ŝx��(�����{�����J�\��O�X~�j�IA���T	�;$��O�����J�C/�U�۪��t���Z���Y�_U���9*Խ�=� Y	S�7��G�3T_$MBw9�w����b<P� W���`��άm�����!z�̥g K*j&Ԁo�������p�toqV���xI�'D��_1Fr9�`�����+?i����&��mS��cP6:�ҳQ�1�|9�J�m#�颸����j~�e�u�"z��E�����HF��^��(�T�T:�8��ߧY�8�OXn�����o��\-:M��RO?����ԟ��*(�%B��EaR�Цn�~��*L�2�B}�m4���Cй��c�%5��!��h?ȁa�M�Q�՝��A_�]b
e���M.t��m��y�%|��
&���wm4�t�~s>�F��T�+�|��E������й]���o��L�4�غ�!�|��ߓ�[�:s�K^�j���W~aɛ�DB�e`�I܇$���K��kƙ<K��d#�Q갰���SĞw�L�>�-,R4Rp�`X����˽)j�-A͟�;E��
UC:b�3������<�9��=� v��Z0�����a�}9��O4.�[z�)�:��Ef�x��jׁw+�����(�d�А���Bc	�A��E|�DT�#-�~;�o��Vn��	a� D����\ƦC��E֩]�f�:���i�de��τ�R܆c�׏Hyh���p�^#P�3��^f;��Gi�����S��!�Ku�2n䖌�F�q*�X�,?��{b2�9ø�f*Bq ��G���5RH1���q.J8k��|b��w|����OEͱ������2 �y�˵p�6��C��?OM�K��Lت��*�4��&5Ȳ�?��e�{��♉�F����0���1�
(��l�e��3�tk�]3dT���T��":ָ�S���5.e U�0 �1S����'׏��}I8h7 E����_���3U�Ð%�N�4Z�ZK-yՄ��t���.,��A��C��5��&U~w��8������~�{���1Q���N
@�{.L�h�����	�-m�1;JXƦ;?.�@.��t�6a|d����5��n�]�z)�������J��چ`��L�����ٴ��k�LT�w ���?���������q��BIK���C�ȱ�hgH�L�g�����w؜���*����7�EK	]�^т��y���J��V�!W ��W���\H�+�D ��Jo���v�i�d؊�H��e/XaX��{�
dny�H!��m����>]-����0�q+
�7w�x��e�b�C��' ��p��W�Uaf=��lo[*9R^"�x�~B�Y��0-�Ƥ�^������ܰS=u��ں�ӶAJ�g���y�Uv����H��t|0�n����#6��+`)�^;���2���Њ�R��^ȫ*G=ѱ�(bW�_Cg���>~�-э��i���zVI�u�So3��1;ѹv�Ll��}̠����ゑ�^|#��tQ���/U"@}`re���*�l��U	�=ү�C*�l���^���m#-��t@A�%l	�#�{O���J�>Y������7
Jm�1}Q#nb��O"���-������X΢�{4����u������"������k�!%	�<���^Ȣ��z Rf�x>�2,Z�%������I�>��=1/��W�%k:�����\��"sQ�u5��K&�VW��J ^���N��vS鐚Z�Ν�C�,�x�0)��Y;����GBtY>�T[/�	�"�֭�9vM���G2H�Ib�Q���L�T/S�ǽ���Vy1�?����c(mH���Rp���\�x;-m+��=�*���#��@��i�l~pɄC��K�oFV�aѶ��URbV�X/�4A��]b�R��.��I��`���b�㽊�㍈�W�;:���z��@��a ��Η@Ӑj���?z2��ƈ���b�RVjxX"?�q83pB������I'�	�5�P�q�U��j o�m[<usG��L��H��kSÇ��dѵ3�.!P	}�&������.�,St����&�da�CY4Y���3Տ\�cB�P0��)S�[�K��!�5I%l�1la�|5�z3D�קYz:���۽����Rߕ�F��Brn�q�Q9����,��|w��������"��N��i�����j���W�t����kw���ɹĜ�Gp��2�R�Q^��2�&^�u�/8�%��9�4�M��S�A���?�wd�f���Dn��HI���~L��X����w'�N�u|E��?�A��d��n�����C�?��f$���f��&�t�x�o���S�]]�x\Iʂ�YJ)���A�`�!�z���0�:��
"��*�8M@�t��ݘK�!�{��S�r��Mڰw�Y�vY�bʺxK{+z��'<��ݽ�A�D��Hg�ټ7+>�o�]��g�2�%&��yz��a'�K�맩����<�>��O��v�#�TW�=NQ�CC��7�X�X����=�)�fgH� ���&w��e�GEa�D�5�}�E`���T��po�;����xCA��>���a��3��\�
- `��}��vejsG�-`��,��gG"Y'?�>��k��2��+���M��$-Cjp������഻��}!�����.N���yU0��C��Wr�pq�=�������`���^��#�o����X&�S��yb�R�1{��0��oE8S��K?D(�,�@��?�y+�\O�k���f�&3[W
�k�˅!.��t���1�X��eP��Τ�ߓ��`ȮK��K�[�Ÿ'֕,i(�-Q��rF�U��o�����3/���C͍�g��	�gc��盶�=1ݩ�+'�8*��l���}X�Rq7��˪-/���3���U����9�}�ۛ��O���n�Er�}w�X\?*��p2�!șk��Źf�:�g��co��^D'������*b"�W�B\�ze����������\�/����,�U����j[�i K"�'Ue<8X*{�$͊7q��O2�Mͪ.G�����Q-��	�I���&=<��я��0�1Ԇhޝe	hЪ�M����&� |>-��y�����s5vC)��y��b� p��J<M`���x7����̥e�B�� n��=w�k*��:�f��R�)����Q�L��M!�@O �PFr�5���-�����&�8�F�;���� /F(��X�6�!.O
o����@�=�<9�!��B%�X��������78����6g.¾a��|��!��:,��G�Q>�m��Xt�!)��C奜4��aw��������?!w��P�Т2&\%��w	�Z�@ȱ��t� b�S#�ۯ^	� �v\�s�Wd\w��SG�Al$����ѕ��1 �өoE�+�23���̭nC{1t�s S[�!���1�w=���^ؙʅ HJ�O��W�޼�o�.�t��y���6��n=mz�5�5f����>��p�}�21�r"���G�����w�ڐ(�,�F��ZeE��,�B❭��
��.x��P���d��چ�$x¢U�~�qŨ���Q`���(X<Aӕ�3�ZF_0BP��o�w�`�zL,oqR�rw�ʹ(!����R%��M������p�	G��l%tPu�W��i����������"��	�#	6����5�+�Z���FT�c���B�ӆ�5�rz�ʅ*�w�I}�Ҙ�M����A*��́*:/�#P�(@Qv��P���j�l���r�Z�G�0�w�_S�x�m3�z��Xd��] Y����b��c
G���M���*�y����F+�����Rv.�%�o�wd�-��`J�w�߳�	��[�5 �:_Y���w����-Đxy��U?h�=�j�����I�����'�vl[�\lxgR� ��*%�N���1�}^J��ɵ��(����jp�?##��}!I:�T���6��K\��74��jo���+�RdN���=�ԧ��@��@J���K|���ӱ���ޠ�4
���{�j]i�;g2-#-u(x�9���3<^�
���$���&�5�V�Y���Pv��⯃
pwW��ޕ��;~{����Ç;�����w������CJ������I{�Y���4�}���آ�*	؂}/~���g�4��x�ŚB�y���2���^�&ƥ�~�Z�E�GӖ�F���q#�����lj�jo�����0m
�kk�!��<�oZҽ�H�qF��E�@���K�J
� FP/�Ή�_a�>��QR��������r6ߛZ�V.(x�,cƨ���Y�ķNa��C�x�^��U7�Q�H��+pw�hC���7m�T�*m������LP��1���ق����`O���J:�wB�X��?�fg��C�ht�Ő:��l{*�}���oW$@��o+��W�5��C���HG4� �=�h��4BT�BB]pH`t�'��v#�a,��@��Q3=��$/Sֶ�'�YӛkIX�mS��V4@��%�V>���D�UP�9���;�5�ŏ�b;�凭"����Y�!b!���bdl �oz�(�Dt^O�U���w��<�z̍�	p�� m9�	�I��R�?�dgqk�-���O�C�~���E�k�E�zd����݃��X�男�(���\&|�-�_B�ę���mSs��#��V�B���~LCNb&�<�3�|�2Ɲ]��_q�f���?BjD'��>u+��o��f�<�8)��S�n"�㯗!	iKC�$#�su�Z��^�q襋�QgKR/�>�X
�^Df!���0��l"���b��G��G�2�aE ���������wZX7�4I�3	͝���a��L��Z0���W�U&�'��%�잞CV�O~�d=)�q!V���r�J�f��X�D���g�"���,E�KO�!ۤ[h�R��5����D%d��][dF�5�ph�氁�a�^�17�PC���;�db.&HBn]\T"��fK�[Z=RTҹݚ(��Ъ��K1��!�������;��@;��'9OCMD<h?�*K!�nAk܅�����iu���]0a9u3@���j�*6NʥT�bc^�fH,��C~#��{�j�n��<����n�Ͱ�* ڣQ��#����7�T'LD�srdӕq�o^L���-��V���%�1��c/oɽ�9s�]��X�����C+���;e7�Hw�2��$�LGI�AJ��K��2��Pw�߱��t�
�{!��rq�ʭ��0�v8�A͉(�rEҗ��8�BtU���s�Xo��GG�ڷ�5��N�a;��	�\�p	9�?�Z �p���C~�ԁҷ���[�bp�]U��w���"�!D����;��$Y0���be;�}�(A]��Q.�JK�Ϝs�+�w	h&^��H���rYCO���Y�f�w\+�Ջ��vw�Q��ˤ�zQ➙D���,��B���LF[���Ӈ���p��.�3�d����C�7�� ��I�����o�����P�\��]�Zx�p��J'���m�#f~��� {ĎU�P�LZ�LmU��7�]QP e�Tఛ�$z`FʓD}ZU
{)Z�Ɨ�OV���|m�D^�f�e�v�E�+OrK_}eW�J�326x"�ʣ���Ыa��R:s�K��ņuuiQ�	�1�U<σ����)��K�?�Y� @F�2{L�?ָ�#VbNZ��iڶί�qρ�Q���ܩ��"�����Y�BJ�S
���`�{��v*�tT�S�>�� �Ov���ۊ�dЉl$i%,x��V�E���u��`��-����WQ(���K�x����[c[�/73��z��8�JI���O7�6H���7"`�I�U����O~���F�����?h�]zgu�Vwo��G�
��ad�y�q4��n�>뵳�x/��OvuA��/���<<2�@��E�(-�Mǃ�&���\ �]�4��V�P6���{$w���+jnS*P�N�>�n�	XD�<�hZ��M���p7)t�r݀�K@\�|O����E��I���|Td��R ��L����,�04ܕ�}2M���q�q�P6��W&���R���6k���-*W���e(���?��2M�y�8��X�6�i9�u,+����$� �pA�;j/�Aq�dJ-�C�Vw�5���HV�.x���^��o���w��f�j�ƅ}��r*@��H�(��&FQ�OQ٫W}�d�nQh���,��3z��t�f�fOVīH9�$R�Tw����c�@�Ro�����&k��)(*a���٘�S�C|�� �|Σ�$�? yT~�80�uZ��79������幦�9N�A�����4ft�׌�ɏ��ʟ6ٓqϐ����� 4�7,ѻ��P�/�A��..�b�)��N�YD�k �ɣs�y�	�"�sP�#zh���)���mcK�O �{���P�VC������*0�$�>���gj`� PB�oY�g�P<�قc�ɭ#�v��yl��p�J�m�$<S�9KωB�;/O��c���ڛ?c8�C���W�a��cC�y�Ż�1��<� �s�!�A��N�S^Q��T�j�a-�qYMF2�P��#7)ߋݛΧ*$d �L�聆�捘63qy{�2$[E;3�rZ%e�(<���lOz��EWu�r������sZt3'�9�U�:)�(Y�Q~M�#��qԙ�I���A܋���1?>��l�*J�%�o8�?�
�h��ᘊ[F�
j��I��)�ٷ�R�1 գE��YI@j���}
�~E<��9�Z6��jG�U��e���t��zZ����C���I��j�v�� &�e#6[���wW�؂ws��.g��7�7P���;�$����zw_�`6TfL���y�#��C]MB�_W,o�dPG��$"C5S�EY�ʯ�$���֘w,/4=r���M� �t�n@�s�p����SeS�{=�ݖ��[���N����>����B���n^����35Q|����I�h���d��Dr�L�0������u�}�/\'�f�b��
(�c�\3p�����>j)���zFp�h�#�-��6��R���, �+O�\�(iV��x}�mQ���H����"u��J|���A�O��� �^���荭]�qP_FV���"�Ʈ�ݼ��� ���'���gxmX��]+I{ q�m.���w�w��������K*�y����8��YӪp�1Y{.��=(JS 9������<�s��n�#^u���U�>������N%W*g�UV NL�jmi�\0U��|���\\Z�K��	��7���y�p��T	G ��� 2N�J��oj�Z�?j��/e(*� ۧ`���o�c`��L����a�Hi�R��n?o�zL�90���@����l)��bE�gOJY�s�5�Ƹg�v8�J�d�r�_)�v��>�.�A��v���F��%ʾ*E�
��Z?��	G��Mb�h����[��旁�b�OG1*3� c�5�����B�c�2A�kFl��(��[絈�e��g>����!��Bmb5nMZ)6�'?�Ģ-B\�{qZR�ݔ�i��~tK��M����-�� '.˲�Jp�^C~@^�E�mN���|�_�E_c^�,�V�=6G;G ����7�K���.S�ҙ6�X��QIT
��/f�[Qf�,�I�P�1[�2>�Ӄ w�p8�{h�4�yxm��W�zٖ�:���E��IGɃ���U��x9N�����������	/Ыv��MW0N��v�u��I��"p]Ahu���;C�A���s���𞞸g	F�M6P�vz' �vm��K���蝫ϒҮ�����	K�;in��)�l��ƅP4* ���-m�,1�t�u���Ys~݋�ջ1S�#�׻�X����Rq�ٙ�s�C�1�P��X���c〄ə���b���P��0�7|�$W�H]�(�θ���V����D���]�3�����B�;��� �2�:5�T�#��K�d���œ����0�s���=��pZˉ��>�m�C����P]�<��W|A3��H������QzHz�e�VtEF��t���P����������r�O��t;�_é���Yx}�r,ٱ�1�,;�����W���&�����̳S&���ܴ�@t1�:_8I�ZיZ�vOv/����WF{z�w�KW��Ѯ�<z�6��7��|<ɳ!V�9@�rN�ͬ�uY#��k��>k�<�����"�/�$�^*���ϰ-@nʏ��:]/�f+���=�F-���k�FE����ȶ�]q>�"Ɇ���(X������,��DU��)R�,KKZ�!�p�
��{h�Q'��]�E�o��׸.��V��߬�����?6�-�g�>��%A�3�f8G�'wzG���'ӯ�z^��W�<�J����6r�w	�^�ey�1��\�ͦ�)�	�u\���c?k<��Q$�v!	��~�2���{��Nx8�����}���D�,v#���=1G(��S���#�o��H��E$`�%���}x�p���q�U^[�����;J�Ϳ|�\��w18q;�˃�v�i!jn�<&a���n�$��\Y� �@MM*�>d%QM�zbF?��,.#/z͞��K�&@x���9��nw�x����R��i���@偊�N����O,x���E�cc��4^���(����p�r�c���K��c�{���[�S�g�5Ԁ��"*,�c�2 c��͓��S��fN���hUyiD��9�킠M�f�8�ת�ӝ�R����rK�7s�&��p�Ă���Z��e�w�=K���"�`H%�h��|����z�!޾gd/>`޷,b���ݩr�ft���Hb�o@���=��f�[z&�z�! �ҝ:�-Вt2�JP�$��d�-��["յWIm��9��X/�L��)����m@�W|{(6�S�ad���/G�f�.A�fbv�� �q���F�ꋊ��Қ�N��`�}�I���y��#�b}P�iٽ7���Nb.�3���2��|W��l�]��O���%��US%����Q Ql���!>'���߸xL�r�k搫��%�R^)�1pn/Z�����C��qBnq�(}�iTh�}5Mdbc��t�Md�M*����C�`G�2��>���hi�X�s��ͿV�9K_��Rg�_��q�&�E�9`Zg�7���cs���-��U�ؠ.*�GԮ�:������d����H�7��G�5�'���#x#�}ۑ��� �=�F�?�W��SqP!r�|���%��	�����'��4������;a��M&�A�:H�+�N5�%"[��tW�o�	�M�1@A�U���"$�nݦ�K�~���P�h́��Tj|�ķX�Ҥ́з��r����)*�#��!j���JU��a�GbesQ��X���e )Ma�tb�6��Ɔ��?�;�
�/� �k�qí�rf��r5�
B��"�s+||b?"���R�t�4���a��y{0K��(�U'��u��M����+y�~��vΚ�� ��2� q�������N�uӔ�C	�jq�(�:%��׎������/��>Ϧ�I�!�`���5U!�<	�����:�P@��;�4j���I���A����w�i!�tǤ쁵��&���@����'���-���<�+����zF ���6��տ;zmT�4Q��Ie�\ݷ}��~"�ï�
��M�����^���o��0n�Bv���}�ҟ��Z��=w�^����m��\2hi�S���FwRz�Ѹv$��z��V�r��idL-ܘy��.���+�?�W-��1\��[��B"��}��v�{��
���N	��w, ��I������Dz6���*�
�>С�^���[��Q��r�ӣ �3_+��Q�\���H �!�����v���%�Z�3
5��������P�IG�cC����*��E��ze�duW�8'�Rm�;a�NK�XO����.�c���kԥ�3<r��K�������&�]![L�/Oɂ�
�QqŘ���������v�P��AI�eK������|r��-zL)��i��+"<=�q����v#�>F�����)��#�53�8J��5<?���C\��;�ʑ�ˬ�2���}��,v�r[c��y��wbX�N�,�wc�粵/`��j
+��Au&	��k>�iM��kM�3������vU�Ƌ��.uC���h���#�Z F3]s��U���vH:?M������;F���C_wSoSӅ��^E�w5�]���B�C!���jd��������Fտ�?Hֽ�Eq�e:b"o~I^�U7��|��!��.��C���U�轼7B���!s7X��U�WK��Mh/�����pI����?�^�E�`˭cw�
�ro�'ܴvb<Y@4Ul������Q���2����Y��q�������1�}��!��eЛv������r �Ey.6�2h��"�kq+_?��o+")j*�"x��=z�� `#�M馲ˮ�K��"�_��KؒX� ��$}_4hb�fX.�d�J.�؇�Q7v*��eڑ�~J��>�_KL�,8ې�"5e�_���
�Wh"����%fK���PM&"3g�y�����"z�)g�q~ҽ�ޒ��$���P�e�s
JT-˘B��i�D��+%�]8�A,
�4�m��[����2��Q��.n�,�T|���ȠbqNPA!/6=��- k�/��m���"���������r�->i  �q�AˋӦ3U���h��\L�_�n��粜�0�~ؑ+�҉�PT��?�%�H�f��5)�[�u�WnfUg-J:x��ɓ��
F�{G&�ˁbhE���QC%�[cQ�%c92� ,�Z���� �&^�
����'���[f����A;�Y�^�/ h_����.���f�s=>��G�@���xk����5�������~F��wlYc��1��Z�^m��Ul��if>��m�e�[n_wRk>!%0���R���b��.[H��%>
�W<�*�IU %�	�R��#�G��V핞���j���Ak���r[�C�;K.y�UC�4A"�ґG�\�./%`ޮ�z�d�p�Hq�|���ga�3�Sv����!и��B�=?�m1�Xe����l%=��'��nMV7S�E�8�r$�8S��g��0Lg��	 k�Y��Ǯ�"D#Щ�MRY��V-�y�8��ࠥ�@'E�k�����8.c�ĭ��v0��k�F8��x�������C����5dR"Hd=J�ȴ�����Y��e[�2��Q�����6U��f��0�C�U�e��@�"[�Q�R���)	�V�~��dL)}:�8f�)au�q��XC>�2�:�k�0��l��6KFm�;�l���{���ƑrL����[Y��Xܸ��e3��9|�b�������<�,q����΂�.==�Ҩ2�B{7��d��.~��Z^�&�k���Lhђ�U�"�:��+?�ݽoUX�-�hd0�#_p,�Fo�Hl�+�R�Tb[SK>B�l�з����%�\���X9�-�OsI{/��G|���K^y7�⥟m3������@1+<{��Yw�����ڃ�x ��p�[OE�O��jT��N8� ��wzH�y�%��y���^�U�y���D3EV�N)
��th���ռK`c�6�yԘb,�K��{�/G;щ�Q�ut6chw�X&1/5kƗ�����N�ۀwo�l��ɋZ������q��,�Q�\��\0�F�D��AaU!��Q����Ą8���Ϲ��X����~��=ԯ	�"�J���{ � ��$��v1� *�	��O܋y�d̙P� �ƅ'�Q������=�(�O��;�L	���;�C�\�Ԋ���""4r%� �GUa���f�60�f(�?���CF���讒]�/�*���.6b�����P�n!��n#���	�IӢ�0�l�fF}`�/�Ͽs1��L���]�X�Q����Lԡ�F\�9k���A�oWz��E��9mXrvÐ�k�{�r���ɫ��Sbu�A!�!����-W�b�1���_���ذ�����#�:J���(`����e��
�i�=
��:����U$?�!	���,���|Ѐ��Y���~�	��i��E�rY)7��n�AO��b�ˇ J���T�9��A��0�����f駫B&ٗC�h.���<�KAe��
6P�9�aY�O�Ä����,-�N�֥lJ��\��z�u6S�XS{fn��w� ec�{��]_��:_`���2*s�B�g1i�r�u�ԅ���D�]�b9ߐf��NGz�U)5T`��p.]l"6���3��@x�O�M*�N��މW�ȍ(�z�Vm�.��<5OS�*�n���-��0���m�~�W�P�s*������;p�����������(��Vd���
��R�q����-�G�m�z�� Z�_�J�d�Wl���z�p�t>�xņ֔D��^�ȏ��<��s��}䀸���41R�^ԍ&Q�	�0����G���@*�9v�{�����N�n;��.gk�gF+�V(p��j�e��,k�G�{�Tm4t�2��9?�:���=��l��^ 3�ޢ!ǼD�㘍�Ҷ�*�Ѥ��H�6\�0��q�����G~�1��hY�oIGO$0��x��C2�X����Nz�7Е�E|��i�)��1Tfq\-�O����7*#(e�ex)ꋧ�-��\�EP'�x����9ˌ'E���t�6�2-!�����i����ݦ�f֡+��l�K����	.�!/����2djgwW��Wλ}Y$���o���R��0��H�η�;dޣ3�;��|V.��@=ߎ$e�.�E����~�^��h��R�� �&Ď}N^Δ0}�w�fͦ*��è�>�:=j�-q(HM��u/FTn�l�]J<�$� 8'��;��#���p����/MY�]��������-���]�.�5*��j9����/�n@�_Jw�eTPFg�a�!@▃`kF�ݷ�a���[Doz2�>����~��irP��j¤ةX�T
� D����6/�̬#e[B���~��rY�0��	Im�j�ɣl�_��ҩ������2ѝ~��L	Ϟ;I�J����L��T��o ���l�!P6y�O��,�K}�6
���'�������S�����Ⱥ"D�Q��j���>�2ԉA��A��eq@���F���,�̒ܐos���E��B��:�|Ȗ�=���@�ϩ�c\Z�y1��Dq�2�(����ܘZ����_��xrqH�s+Xc�ê���G�z�&T�o%2b�Am�2�.un{��:�b�{j���MԼPO�V�I��
ܩC_��4��|��i�����x�i�I(q2}����P%;�����/��������>Tk �6�G�+�~؄2�a��"�������J����B���9{n� UИRu*+��ȃ�@+�SR�H!Ζ�{��i3s���cu )�D���<1�&�pr�NZ��C�jftAj*2��4B<�p���
*��Pz��9�0��?�����x�L��CD������6t��.�dp��o�$�I+{u�΅�=u��S`��*%����\w����/�c���w�=���rT�5�tC'Z P�T��6+�ku�%{u�D'%��!�ۤ�@U�X�Lu?�
8$�C#J�)�w@�А5|�m$΁���z���ز���o��1s	�`�nh�� �J�ˮ�Yb��X��5�u�r.���;����3�Ē��-J�.s�NԄ���D�����1(��gj������xt�d̳U��s�z<:��Ljy�z���EQIz	��m ǃ��
6_9�wI�����r"q��9��<�T����sTq��h�U�Ҧ�=��U�}�3���@5Xˑ֯Zn������£��2wn"�L�obѷ��� �:�ϥ�q����[��7��9��2ZE뮔'�]���{N~x��X��uE�k�:�۫^�">�a|2��n-wiX�G~g���揹�mC��V�uAGJr*x�:�{��ۆ�S��w8��(U��~
'�ۂ��rM��P���cع�)8��֎�]F�M��z�c!zb���f!���Nd��x�J�}x�D���y笙��6H$�%wZ��[%�����-��z���`�AW}�"�;C��H��bfO�DP�����z��*�,�C�>,q���m��&yO�#�O�ʔ�@�@j}��+e�"���u΋����9�>�@���B���? r�7d�m�E�/���Ƙ<����>a�6��^]%5�9������+�̳�ua��	� X��n$m���c�,D���r��S��NH��I�Va���m�t��?�?�|M�9$>�U��҂G�UX��`�Cyw�=y��}�j�T�N�n	Lr*������������yGŮf�}V}팧��C�V�{�O��.������o�
.2�7Y񩚂������Gp��1��eZJo�~��!�x�
���Rj�v����$���
��ԉ�~;�HH��Ax_��&�ڭ�����c�ŗ�<,-��T�c�-�ex����+%_�)�v�q<\�3�g���j�����i�àC�~�xx����ƣ(���S��0qL8�p|��#׫M̬J1փ�x$#��҈�(��M�k���D,��m�����ya�;9~��й��&+�04���k ����c�9��	���c��M�ؖޜ���e�,T3֨��j���rgY��
ڇs���95D�Y��I�(/�l	���fB�~~���~O+���s/���o�:�%�mm���O���.��@u�7��?=�F��*�mWD��[�p���Jj�Cm�D�O��g�mh��؃đa��_��7�1ϟM�DN*8��-���N����gGR5�Bٍ�E�	�c!3�AKg�C#'�vP�����u(��imIۃT�����a~q���J�ӿ$���Z&O*�m������02���S�=��pv"UR`��Z��PR�tJ"_й�<)ݜ����7"�L��ɐa
�i��S�� )�o�`q���U��r��zT���;r_/�)a�NBb�#.}g��q��Z��P����c�3���ES�X�����*p}/��%��G���SL1ic~��Ū��Ua�n�7��Gg���I�/{�N|ky�ß��-��_�]��Ls�}/Q!���	S1C�9CW�CiY�M4�����V���7���2�����:��K�U]��u��Y��/sB�X�M\m*J���͙�f6>��0�u��#%�	?f?o,c�%�*#����5�9n:�s�J��˳dg;|?�d�V�?c�q����}+�I��,���ch�H��M�,	]^~M�#z��O��e��|w7b|>'���ʄ��>b�M2P������<⒣eo��
�:=t]�V���^
�~��zյOr���6�%����g�o�Qs̉�]�n[�D�d�]��Z�ir�ݮ��lv�)3,�dx��>��gx�����h�;�V�BK���!��Վ 'V������U�s;!$�3O��3��#K�Hd܇�-D�.��vt_�Qz-���������6�V[K�eDԔ�P`T�g|��JI��D��0J�!ɴ�p�q�j���d�� ��S�Շ���@�b����ݖ���)L�kU���*�W����6T���"໷n���Z�'���-���\�ϼHx�/�/cx
�A��-���Bsh
Cy���Y��}�eMw&0�C������3���C���'l����3FJ˟#��^G(�t$�hI\&<!�B�t�9[?O���Xy�e,2cѻ����5��������3̄w��m�c{�/����D�4i`�h>�����"� 7ȍ�i�ӜV$8@7�(�������J�3��D��ۦ8�q2oʩ�e�ab���f@�\�|���-�oJ���l��w�
�^�)�s�10�=ZL��"*��._ŗ�u��O�Ra�8��|����t�7!F���я�%�蔁e��^"�)�M�W�=XŰ�QNN��@ض�z�����=�Q6uQ��p�w}�VŨ��|:�/����ڊ]���2>�P-�zD�T!�������%���@���W��fD ��N��AUϝ��6�?DEJ[@lc����~��e��3�x���ѽ�=��%v�$���E�qd~P`�~��&"��{�O�t3z�8��$�ՙ�����2%��� �hy�	Zd|^��Ik�Q����B	�&#Uw�6�C
���D'Qi$X�D�q	�d��\�p��2פ��w)a��j�qi��B�[�w�Ӗn$i~a����R��{�Z�:r$c�^Q4�ͺ�i�ع֦�h�E�v�A>Ȱ%`'�c���V������U���(��z��,��4�"�˅w~�02����#Q��S��1|��M��m��uo#sVVi�<�y�R9�7� �/љMy��>oM5
ɷ6IJGꦹ:���@� ����-p��.�_X���B���A�Q��q��(��1ۉ�qmh��G�Bq�Ր�w�n�(4�9�㦃fpXf!��UHR������1���y,q�X��F���k�������ݍ��|�fC���"�t'���D:n��h��{h���NNq�;��c�̑�=B��sp���J���� (�ï���C��4��W��q�[J�<�㙻������:���m	x?�|&�ǫAm���ڴ����@`㏂EP�}U�اƴXuY\z=縴ڱ��+��Sf=�A,�w9�F�TbKp�>񇦻^�Y�n���%k�'��d^��c-�s��ׇqX,�4)��z�����ʭ�iM���0L�[���1�9ZC��[��ι�E�9D�M�"&���D�}j*�Ne����oze6��ݾ��>d�fG��=M�B�w_��<j�i���17ir�5�fa�^	���A+��AT��)���-��xCn�<Z� X��J+
&(b�X܇;߾pHM������Đuz ����J�aK 'iN�7�h�����w�t�|=��6�f��R@��t��3��D$,�j�Ywѻ�'��n�!��瀚�3��P08�:������9*�@zg��X���Ņɤ�|xa��;�J�,]w"�9C,��r��+�s`R��[d\�%�Ie/���u��M�^֬��1����>�ϝU;BV-��N|6�j�j�����.FpA�Og�����|�����'	p�
�M�ߡb����@���Me3Y�c�d!�Y�̉^1�.��[�[�?���_`y���j�`Uu�3Lm�P�w��R��ܱ�b��},|D��/�^;X�$)��,�A�\����6��{f�>�IW�&L�]d@��/�j�Z�d~�q��}<���f1�_܂S��E��i�GVY{%7M �U�T����v8���J@�R�s��P!8�jRx�S�D30�3������ �P_u6��iB���06�.��&�l;��qX�1�*p�W��&U���j�D����Q�TL�]eK���|�=d�3i���O��!�-,^227�N婌�DO/N�����P�ëƭ�'�0r�����n@TrQ�Q�,)�Ԣ�U/)��rB��f<����9V�.w�p)Լ�
Z��;^#�0�R$]�g�Q�e1<bu�� � u�Զ?�Z>K�����몪 7��X�=�Bf�dU�.1�n>1����![�QEe�*�엓�ҡ�q���^�@��ObMgX7�v�
3W@��M�	g��g4�অ�R������de��A-�5#l�E'��Zp�#ѷ��n�>=u#��C,�ί<M�[Xj1�6I�����HiDz�{�0BMo8�D&eB�Ȍ���n�)z7�<L�^oP$�9�A{|�V�8М�i��;��Y� �l�p��L�\�5�T�O�ƗƤO	�j��!��H��z ��y{�͢���h�g���+K��]d��D���Rh9�3�� �:�S3(>;����qA&�g�>#	�,e��DL�\x���_|�P��[W���Q,�P�,dt'������W<�<��U�ċ	l^�}�_IWȕ��?���d�uY&��9��~��t���f�sȕm�>����j1�ߨ�N�H+Ry"o�'���-�����'Q��>2��k!у8�,�Y��H8Y$�W�p�}רr����q�P���_��qƋ6�����R(&}K�Z�&˦5;~ׄ`�*�5������M�\z=8����n �M�I����ʰW�`ް:�z�d�a�6i#�8_��� ��{��$Ϻ�,kbԆ�� bl"q����W�$����v��Ѭ���!JS��)������Z�7\N� ���L���[�tt�s�"�HqK��F���c��4�����4w�n5p%�D��Q���R������힪.X�De���?�([*���Aߋ�m�m�u��o���&�_�@�\�)���|��ۈ��*f���Q8�@i��K7���K97��t/�'�m��ۻ�0Q�p�(�q�B�#��P�\Ak;�St�z�汁�<A�DHs��c��i���:ν��jݎ4C���*9�'�g�ԋ���H��e��Ї�����㔟��(��v��SC�MSͽU�g��#%\�]�+��38M�^k�@���٪F�~�;~��7�F���M��Kh�:46dzJ��P6i.m�]�����Η�h��;��Ԇ�a>���V���e�W\�0k�J]?��u��lg�B�j�����%:S�uJsYy<��+�$�w���m�: *%/��L��w����2t�	]S�ѐm����y���0#���?vB
Di9�8���&2�]��F�[�<�J��?��Eq���:��K�^����2���_F�<=�y�7Ƒ8��^|�Q�hQKAmQ�I�qг׋<4澶�#8���T�0��mb<
��d�n��Ց^�;PWp��6�M���A���x �L��)�����y�u�����1BAP���9�� �j�� TLE1�豹�W}�l^rz�iR���{rӻu�KG�����s:��PA�I�N��}��k����D��x^�)��4�u��T�۔(lA�ߍ��ȹZ$_� h�w��znXC����C
S+V�}65�e�[N�t���е3߹�#_��í hԮ�3m�Q����q��ϊ���{�q\'5��)VbPC�K�W~֮e��lp����>��C�fN/�hw�@]�Ѯ^ze%0����F�$?Eȳ�=��%30��{.KF1���T\�2�N=�>ǽ���"0k]�(,G�Y{��A�Fn[���h%�!�3�����/ͳ�|4�������!�ݺ�K�!~�o�5o:S�.�9<a;2��Zԝ�����b>,�j�?Le�'��P�"���:!��c'�]�$�
��e� h��(�F�(�l��Ĉft�f�ldw��[�uiă!9ֻ�'&��v�]�{��$U�������r[>@I�}JBg�8����0��"B�ᑦ R���
��O�}s��[��J����/���f�p+ֆ
ͻ�����@m���ҡ��߁�gRѰIm%�2>��s�d�&\�/�����}|�C(�Ӽ�7C�7/8*�TlR$<���~G�^:VU��tҥ�����^�!�K��*������������UW��B��ȧw�蟍N���/>C`H;�=S]�`7��):W��o��Z����]5���4}�R)T����k����&���wp(�ա�Ȋ��6�<�T�־�r~��o.ɛ�� 
RV�?�mw�����K٠˫�dvvs�(�"�]p��"�YQ7$��:���v0�\�$Kӷ����IఢYmOr�8�C
wa:7.�p�Ñ:;��p0�Ր`F/a��yFNz2�+�LWBǥKb$Z���gc��m<:�K�M��l>�DӅ�!	P���=���m��+&����B�Ti�\�%z�hX,���)��>�ʻ\�u����=�?1}Ze���O�mX��~�
ϬW�	�ûڹ�_�|�9�U�T϶����Pձ�}��R��_��|��Dtٓ!ki5@�_�T��\~q.g��]�/)A����c��D�<��A_!��
�e�n�n��v���j�%���^%L��i�-�I.�Ӏ���&ZOf�RM�l�- �D�`��Jפu�Z�v$�.k��:� �B�/k)� Au~���-��)����·C��y�:Q㝱����i����
&wz3��؍`NW���v��E�W�T����F����G¤P~܉$D]���[�1�Dk��XԖ�%mz�h�Jɜpv�[�Dz���$�.n`Mӛ����L�Jq��>L M�7�T�_[�̐9CXyebwB�2�c��?( ��I~M����"[r�C�~�6��b1YIA���V-&%4@������3h�Z�"`/Q��$m�Շ��fP3��UP"|r1A�����.�x��q O�|yX���Jy�V��#����pW���¸��?���F<�!+#y��$Gy�?$�)GK�-1S��##�̓c����E.󗜽|]?[�Fkss�Zgz)*d�+�JOl.�z0��Vᾤ^�~�G��NRT�:l~֣�_�}Is�����Yh���_w��AW�6)v��{�w�u��>��&����$�N�+%�?�7yU���c���B䁒 I���V����)��gE����:�fHTdV��D��e��>��gT�-��%�"W�L��|e��L�����]��1�#�}QB`��X�Q�a?�0�-��w��8Գ��_@�����=~�+�c�]r3�AO��v��2Z����Ǡ67���۩�4��D���Cr��z�T5X�Z��u��%��'���_�H� ;�c^薰�3pP��x�\� ���tX[�(�H�¿Z�C`?˧��}[a��[�2��T�S��)A�.�*�.gZ�AF�r�}}j�HE���x4s�yU���=3�6ES�]@��8ԉ�C����&�X��׎��g�!N���h4�e��O��r82j��ysVUMf<a��u�nJ6U�m_G�#IwH���!g�{f׿�v-G;�2ś�Pդ�dNG��U�6{ g��b�[N]&�J��ݻVZ�m����H`�7l��xl����L�%^Q��\\���&�}����5��+��\��d �3X�!�N x^�|����0?r�n�5��-�U{�����Sư�vc��oߠb\�N��)ɮ�kp���~X��A���L��@k5i�d�,8��>}����>�2=cLX���6� (��@��G��H�5f����W���+b0����%ժ�AZSU/4w1��E+����e���Q�iL��at@���P��۪��C'��	e�F��@SIx_Y1ª���e%�s�Ԑ#w�0j���o�rK�* C�q*(2'�?fv4�!�ò�e��X��|�8�w+�R-�-�-�g�&U�un��t�4����`�_�(��|�	�"�.^��·yyցw���Z[�*g9�zj���4�%���Uo��	'��Z��G-2ڄ�MvX*�T�5��9뻿�t�XC�Tk?�y�}k�G�o7�AѦE�$�0/�W��0f� A���C2gb�IQaHL��*�����
#��-`1�/�rqR�&6�C�!��șI@?L%��~ί<�`T
��>��yS�! ,��`A�2��b��%������-�n��3�@gn1���5��rY���]��5ʥs7̫+�8�w��E䴫�^�
�@�/Ss��=�!âc�$`��A��Z��
˺C���š� I-ј����3� /����"���I��T��`V�ϤX&�����4�N8�����$�1v.���b��X��x6_c�iT:�����2�n���K�u喧W�Ӌk�(+�� }w��`�,F����z-��r��:M�oU"�D,��+��@}h�`�����y�/~�F|}�%���&�k�6��M���/�jd��0c����1n28S��;"��v��f�J���v����6����զ��Teݾ�:��<�7g��6 ������h�"��$4�ՙűl\��@1�!8�H�8�"�	�PK�<Ct�Я"g������i�7�8��7�!Jj�����G�i_�Y���@�}���n?�#>B���ұjS�-��bt�~�<�m���O6r�!�Co�oq`A>ViB[N���'�^��lτ����Q4��˽4~�g�ⰠUp&G����]3��W+G�H��VN�b�&����&�7���<m�h�P:�s%X�g�"M)N��λ�%`�I�a����;*�p`�y��x\z+�4o�*�@n\��PW���1�)�����KT��Hy��hh�Ğ����!˙��.��.r�
�/߱[�j,Ѷc��L�i�Ř�C�����iC��BxFz���|�U�9�"\ڜ=��1��ep��`	���V�`Ѡ�h�}a1�˛mي>3Uhu+]Qn
�.������b��D�0O��Q�%k��K��ǟ�63_M���$>7*��[\טk�'c�:��6/������Y'{�)��A�g e��u�|G6	���ہ�82Ec��Ǫ��`�D]����e�>�+��ݏ�xx��o�ø�d�f�9]�*��h)Np���]����}���O�G�-,�����3e;��GL��_[R�4!
����U���ZDS�������F�
�r�0UMm�;�ɀ�9���w�5B��s5$�����+S_4�������Z(Y�b�`Aö'���[�R����Q -���^��D�7�����x�Ŷ2�&����,G�ǳ�>]Y(�J��!agQ���5����7Si��� ���"xiv��������w(�)z��������"�FN�pU�6s�b1'f� �hn̥6�a[�h��$^?�oD��������'���A ��}���y�0���:@�� �,��������g��.�z߾>t�"�)3CLt��<S���5m���fx9S(�xV,'��נnB8�(,�!�K�9�V����/��]y�>Bx�u^!� �y���%�Xa���J��n��q����#�l�;��d7���4�����MU�~u�SO�FVK�oȋ��@�W�6&��L��I��%�α��iUZ%���2�W��=מ]�	�r�v����9�T��,h���d/�*�4�
�J�x���G���]��U����� ��	�'8��RE=�4�\�����JnY;�o��+�Yc0�����m̡��ʉy�jnʥXƃy���h��X�y;淵N�D���5Q!R
��BG��~��|�����J�H3�uB~K=�(�F��"?�E�Y�ڜP]^Y
���@J+�Z�P�sy4N�P��c�8ҡ�E���E��`��5,�#{XRi��gO*�߈/L1f���8���;�>BĚ׺�#@�؄�&��}/�uA�H���Y1RQd�f~�j��oM�4��6U�is���I��"��a�Sv��{��w �1���h��?*�1Gi�/{lM��.u\{�%+Ҝ���Ґc���.j�S=S�yЅN��M��k��3������)��b�b?���Q�x���)Pyh֑�.�G[v禬7I��|�o�og�,7-�C��B1@�	ͤaM��VS�n%�l�~OTOOY4���s��n 4l+�� ��R"�%Y��cf�$�Eܕ����?�,1�Q�l�,�ܠ��2��c��
�Ԫs.��!��V�5�0N�kD���^��4T��ڃ��\-z�	$������Z���)���.��Y~f��KY���[���+�\�?�'�4�J=�tż#�j���ٌ�j�Y�An�O(��ٴT�ǡ�j��N��o��={�M�F^b2��l������%�;r�{ޟ_A���r��BӮ`��K�X"�9f:�r�og_��FӋ���	;���F��i*IT���蠒�!gGs8N�L��� �ݝV��x��0�}$��0��pR���	J@ʒ&$;O�"�o��W�&�{���ʻ�zq�B� �G��ɓc)��T*{>���9�����g�ᄶFcȁ	=ݠ�R#�A6�z��S�5���#r!���������8�3H���J�:���<���̌�ױ�^�#��"��h��"�P�`8�����iW��f�I�CS�: ߰q��;T+_�Nsj���N�XW�NFcΓ�U��,��&Y��5c�L�$G�yʁ�� ��<l��Q*����+$a�������v�U��>��J��3 HmcM+A��m����1x�u���\	�x�3�Xĕ3�IA�kL��!��m�����{r���ߟ5L�W);��X��2\9>1l��C�h�����Q�c~?�=v݃%���5�u���Њ�qQ`6^���~L�*~8 K�	���6Coݮ:�a�x4�:�?�n�P~���^��ʂ/�Ϟ!v�~����Iq�s���f����a	�"�h�$h�����de1>a<吺O�F��6Vx^�4���e��uN�^��G.������$�Dܟ!�d���Y����9�8�?�Jkh���|�t�&6득����M�냡\I�0���Jԣ���!=��Q���Sp�~��j�~�����0@��v2%"�"o�������a/>?����0k���>�m��ފZȷ���nÀ�T�llp�Z7wPY�^Jb'.ǓY��6 Kx�K�E[����)64�|�+��>"w�IK �?�����`���Z�,�6m���k���%?ڽS<ن����)
;q�Ȳ�Anof|�((�۟:	FY��T�9hĽ`ʤU�3+����e{���_�[+�t]"������ٮ�^S���l7]!&�Bf�#�Qc�>�(=�>Js��$��ELh�7�s����|�*�B'��;�w�M�wr��D=n�..:$\�!Wn���Q#�d	��+r2g� ˴�ֵ��+Pru��1��섶�w�n*|`?����%/,��Mĸ����%��fu�w��!���Ԧ����z)���)Z �?i��N3�l��>��I���Tb��}�;UfhX2�����v�ǀX����Y�� YYcI�FM�Ձ��Jk����O�����gq���ݧޣ���1h6��0f�t��y�]�@�b�[��=��v�6�lP[}#j;DZ�C�������>�_���0fA5���)}"EM�9������O�����ˊ&�Mst�ğ���F�w�����eS6��u�e�S��a��|�P��9DØ�K�@�)�1�`�|�wLa��Ť'�m�Ԕ�V��wd|�v�lϾ���?[�Q��+�8���E��vE���)�ٍ�9�e04���X�a�V��}��?O��^��m������'����ʆ�5�����z �������VSv�"��Z�ݣ�C%:[sj7 }�'�E�݌��A���b
{e�+d�Ƚ�s�rމ��*����6���nK�z���lz8���]hZ�˪Oײ��%��J���q�r2w;؞uy/�ݲ�q�$��i_���Գ��ͻm��ۖ�|W4�Y����`B���e�-Z@��= �a@�¸�FK}�����ā�`
�T��ܜ��򶀱�[��Y�O��-6l��V�a������*yJ�zB���e��f����>����=J�S�������}��!�g%��u><8k#�P�G9E�$	���Ԉ
�v�J�r�B��d.|����&����:e���*�"-pPH� R=����{�5M� ���Rx�Zb���B���h"�z/dc��<)��6�m�����k��Y�D9���r!%� ��"���|!V�M�Ѧ��b�S{���[�O��|)��N��U%��*ǹ����\t6,3��U� ��E�C8����@h�1�rW��ڈ�R_ �S:eg<�F#w�T�L�@=���-gM���Hq��ROb_��g%�z�O	��P�V�Ҩ!ސ<ns{4�p��)J?��8�+Dː�+��"$�?��^�
���3�8ܒ��pj %��o�͒3�C�Cg���B�H�+�������.&��)h��S�/Tx���3�d��_�ơ���Z�h⥃��M�UT��U��/��Z�pȸ�ar]&��ǵlZ��}+rXzL��U����L���"��j��*���R��wx�Zz����p1WXi�\>�g[��/��紦��mbV��y�C�) P�r(u�;����)<���A�B�����ep�K�u��v�j��Elg�dힹ�T��(�#V�q��}��`��E�ؘ��z6���[��@&1$��e JH)�ͱ�R^�A=�Y2;H�R��D�ْ��9C(ЯF��_��x�]��Y��t߫{�
?s>��9����NI��������$oatk�uӧѯ����F�4 n���^c4	*����j����؛V!�w�2���,@��'X�= �_5��=*dbL�����+�B�{�V��}�0g�I�9�⭔LQ�W���$x�2V�`���q�HO�.#8�?���}lyj~��<�0=�c�+�*�8'�
9~����S�z9�g(�
 ������d;�N�T�U����&����'Q?�4��jT����K�`��S�+@���)e��[IfR[��9��[�])�{Ƒ 0���q3���Œ?�ʞ�>bB�D6��I����ֺ粭�Se��U�\VH�2Z��ߤ��K�d�h��p����怇�ͩ!N:�~HMa	��n~�'�d3���z��G�2�fk ����tG�Z�>(Rh���O�.����]�/]o����c����
ͬ�2��5��O��ā�*e��[���Key����zj9 �j' �d��+��/��x����Y˱[jv���;r�0A���6&z�e+�D-����`.쩡�D0�t*̟!��������j�R��E��u�?z)��ܞi�G�^1�I�;��a]�K�ZRNR�A���`NS	̗V�dP��!�~�T1&uZ8^�;�y\4�_q�yes���A�D�5�e
�'u�7r#�W �]E����u�/'�� �*�@���=�sB�󓝕K�$��k�FI︾ѽְ�K��<tD!�<\KG��vB�vjF"~e1��.�;��s���%�ej�0�	��'�B�B�(8�Oh�
���S���9qq-�Q��9���E��	�G3�ⱡ~4����7���[_���r�M�s��1����cCvo��&�a+�s���aBrt8�~2ҕ���K�1��1��`4�g�-(������O(�&����/�*�6�s����OJfK�|�tЛ��a�����MH���Y�ńbn��+��%j*���0D�|HJm�W�5��������c~U����!]��#�':9����	�s?�82��������)z����9�h?�K�3Brg��B/s���:5V�O�̤��tT8�8�GL�7�D��� �K:فl\��������rӆ�9{�[�s]��$s��u6L	�4���$7�9V�]�$f��]l*�m��x�Q2���p"2����j)����I;�<خmn����Ce9���:m�c�I/'(ٺ�%��S�Nތ�dk�g�+N��m�k��:�j��+��E)3��
M{؜HCL�9�L0�%��@D��c��|�pX��/۪4��24ڣ=��4%&l;�1�E��n��w9�<��#��c�-�l����WИ���"= ���xn`�?�Ax�� ���B�&������/|L��Q�sk[��8��ʙ����,���E++"Wk�LD+_����:�LF�x�-=�"��n�*oV��T>��ϐv�U� �h-p�mʽ�?;-����awX�����a���#��G�I$U$��q�D		l���x#�xK�H�<�Z*�G�Æwo7�H�i�4��ᙌK���ޜ������ڑ?O��(~���q�;nI���y�r�����7}|��u��]!���`�3D�b�S�UZU |[0������; �2�������_�6`���\���Da�J^-�k���74������D���JI��4k���<
�yK��0��]��-i(��WR%R��Y����TRk�N�����,S����)�!����N�c�{�L�-z�)�H#^w�fn�?(��vMw���s��:������%0@u�
Abr���r9���;�;?ǒ��yⰦ�"ɦ�t8*b�+�Bo�Tf>S��+�_zœщ�,��q�/' -��O��߭L��[0�`%���4+��J��𴨷���ϡ��|���8���|��jI���w` RR�fo�G�:�i����l^�F9C 4���I'�͕-�7B~���I�[0�
�9���q?�~4��9�����]R%�#;!4 zd95f�R�N�&�-dn2(��(���[A�k¼�~	qH��r���d���p��2͓?{>ܯ��	ɎH��n��z��a�N<���8`t�;�~�@��P�M=�f?�jc��L���=7z��1���æ���}>}p������H�����yk����Ei�[�����֖4�r̯�t?����DA�0(ɥ�5v��4�g�
�����;s�x������B��rZkY�e����':��%/L8g�a� �W�ٝ��f;���ߐS�yn�n�ׅ��snl�V�A�Bȋ�.'|s�����:�<Ny$r_%��zbk���0zG�v=aq+3��m$g,���4��l�pZ�8 ��k��<����U��o�u�^DQ�Q�"Q��t{�3x����N#x�xv��,W���{QV��l��[D� 9���]�@)		AM� ����i���4��RL��z2�/Fq^�5��XcU?� p��q9?�F@�� ��u�!c��r� 6@�53o�J����RD4���+'�τiM\��QeK�$?a½�l輜��U �j���sm6R��j�<C�j�ىӾ�"e4no��a_��w$�h�&>"��u�����I�;»�D�X�&�6B�"j>�����uuVfA�!�p�PvkU����(qp�:o�ˍxU�Mv��.��yu��YSe�W_�D�'me��pZ�+�d�����HV[Wu�n�^V�Yl;���y\�!L-DQDP��J��6{ܶ�h�Esox<;�՘�&�F����B$��	6x�\�X^#xqv��#(ba�|=y]�N������U�V��L랞9!��H�[o��Ke��((!�!�NX]R��Ҷ,�G��d�&qnp���b�PE�I\:U�3�?X�L�݌#�U
[�/� �	t��������`�O|�|~�	�ìk�6�H5����:ZO�}
m)Z�֢~Y �̫�p:Q(���k��Z�߷��Ξ��d{sN�]������?���S5Fs|5�"���'�U_(��} T�vq�M��M��	�.v5m��fձS<9Y��^[�P����1lE�!ɸܮ��?�xh�^!^]��n_���e3G�%��e(���PgI<N��c���τ��A$!uB	�~��P��w%l�,�7y����y���<����H �p��(�:����Htx����CQ�T����f��Z�`�����CyP�p�%�S#��'3�ǌ��$H�p�iO���,eBW֜�s�$�A��>�D��Nx/u!\ސ6�J�XB��Wcڨ�!DJ�}����kO�C���C}���M>?LeB�����f�\ڏ���
(|u�������NO��Jk�w��=f�MI�ȫi��Ӥp�S�~�]���P$T����J
WT�X�5f�ύ�몆��UF�!5������Y�	֘��1����N�+�>�[OO��y���wB$W4�c����#����W*�ф��r��X4l�z�SPr�a{<Y�vQl���T��vhf����i�8���������
���+IZ_u:�/c��L�h�f������b�9=��nHB�"�#e��\�1j�1�1:V�+i�)�"�P( ����}�8h���ϣG�16Pc\�Y���,���)��.}b���;�u��Q�/�p���Lr���oa�������p��/���,�q.����ޣ;��ڗ-_�hZ�\�A��/mo~6����(��0b9���_��
l!�Д��H���k��=�)���j�}?1N3X� -�,hښ*��Y��ԛ�7���߉��_;��D=P�e�W�#Y�h��D�k����a+|4K�Q�O{���L ]p��k�Φ��ɀVM��YxVa��GO *~�*f�A�������3�b\�~<��/f�{�F���Eg��0mx����G?�4��P��5��Ϯ�SPՐ`?/����]�{���v�.���$Zߤ�^�ˣ��=�OT�&h���� ��~{���u�O9�v����ҍ� l�	�;��])�aǜ�����:-��QɮK��\L��#yͪ>�qS��Y�"��_��=�}��f^�@i�]W��/(>#b�{Rp6�]�!|�Xy�bU^ A� �xR��I�=�B�ʟSk�����⽪7��!q6���ԗ�o��i�
�@/z���	۷fwS ��v{�c��?W�=�L+	ze=�ڻ^���r��Q�V��4��}�Y��x��t 
`v��"W�0�x��_� L��w�bzQS�Og��JY�"B��H������������%2��0229��8�.����7D��>�ۂm����}@8��h��M{�H�Y�(�Ō���@fN��8"זp�}0�"R���|ǲ�z�6���b�9����%��&���5�7m�F�(�9�TS�Ni�<�[����&_O(�:Ik�isЌ���1�Er�  �3���l�$5�������)�0�ܚ��xzvl�(a�xH<g��	��9�-���I��l���M��������1�m��x�͔�MS�������/�Z��s��W'M#��G�I+X(�)5�;Y���P���̼�pԛ���VS\~�V���S�K&ue�ް��ev�Ǆ(&���)BJ��-�>y�dmg�Q�̕#ݚ>KM4fQ�Ht�Al�c��Wc��VL��V�Ha7�a��t�E�$?�3�L�VA����Y,6����*ݥ��\tAM�qiB�jj@c�V��f��AD�L�mfK���>!^��h��hP�Ib��\��36P�k.Z�u|�ŝ�v�-@��l��!?��3?��Mg��Q��ՠ%���o�r�7�勂n��P�
��Bs��:�ښP/Qs����h�0�ԷY��<�<r�0.���U�.��~�er�����C:�}�i���7��ˈo��d�	)@�B6���?
ן_����|���2�5bh�
�z��'ӴV����2٘"O���X�_Q�Y�г-�6���!J����^��Y��2%MǪ!y~�|_�}͖�����ʒp��m��M.�6�v�~�5�c�B�w��T�nv?8sNE��9?�w�9[fO���t��Φ�U�}�T�r�_�-�\;OX�hB��u}K�X�@���8�v��x�H���n��"�yW[�v؍a�Y�,^���I���<��m�w��ne�oha�텏
)�Jv&Ǜ��u����y��w�Y~(g0U7��ס:��=:�ԑe��ު��K��6�:��v�x�m�.��X3AșE�V!���qn��fP8�%/��֟*p}I-�Ů��79��	��,>X|�d�L��Q�����Оa����i� Fd�e 6�ʇ�3l�'�[2 e�RJH���+��c���]Z��A�U�u�n�t�qF4���v;h!�7�@^){�W�A����R�$����A����4����"g�6���G���d��C�t����f8I"(𞟪�����5�x8��m� )�jMuןo;Gݮ�1G��dT�
�.8�f�N��a�&u wT��T���I l���g#�[$iD�8�J���Vwn�#X����f�&8RR_��D>����-B����C" ��7��a���vf�V4�(D�Jط��:�_�wM������LA��L8�6P���N [��B#��x�����hl���D%H�+�W��+�\U��M8��A��ѫ���1�><w�"m��|�(ZY�,f�ϟ>M�����F�n\��^�D��:��۴�Mj|���� ��FEG�G��k8�a�
q�	�(��p�����@����έ������FN�)yS�h*Q����js���:Ġ�&�����"$\��
���ݮ--�:m��'���}I�6Y6��L�T�b��Dï$���w���,�	yF��)��c�����x�}n�ϊ�y;^���R���GQ��PXQl���YH�7�0���o�\=uU�o�Vs)7˔*Hg�6(b��^tp��
b~ppz��'�}�bE@v��"D�Ux`E�=YV"��[#�����P�OtE0���36r���s,V��^��ש��"h���>צj:)bW8���4�1�R�O�t��B9�?��g%9���+N檌�k����5tٟS��l-�@�_����Y�o,HK�,�>��̏�縿�5��aY��'j���W�X�Ťj)2(�_'H幨	���2�H��b	��4gL�3����+��W����!��`_���l���K�9����1OШnV�� {�c08̞�p2Y+
Ғ���}.�e��$y��y�P\:�zR�I�ɬvZ�x㔡�tc��D��J���g��0
@J�"N��Bz[��\V�ks�i�6�G�%�	ʟ]1ӻDO{��4��	Q����C'ɗ���c��>�HB*�#���� �Khd��l�����	#4���X,a*8�L:$g����:��G$È��\��`4��:��܎�ebq�)yym�l�-�1�����1�9z�=�N����Aړ6ڠW��BOՑ������N1P�W]����E>f�L.��Z$�����n�QYH�
�4�sd(��w�41�;�'�ssp%��u�� �R��20���/8^4l1���')v�U��8$@�N���1阗b��r �,��6�F�3�Dd��<����;Ͱ�Ɍ�i|? H���^/����⇈)�f:1Fh]ww6���O��n>�:͛-z��9�OH��Vqu�(i-3J�]���5�nF���mX��#�3r�Fu�%�⭬&�wK�h�<�Nɻ6wP�,eW�����e�n��#C�fW����
	�5��Y�`���$�䑊q���C�v1���~���:�AWnO��+����/��v|۶�h���VV��B�9��}��a��(p@��+����Z*��s���Gɫ�� W� 4����`�>E�<��i��W�!z� �l�m�d������Gc���ćT%�]����,+���,ո��Gg��7��o����'Ӑ�&���.����XN���k��1���|;�N��4�Tŭc'�C��U�������{K�Z�#x�> qQh��ǈ��#��H�J���q ��S��ʻ�  �%�z��!o:��Č[��*?쭜��a�E��^	Lni���i����(@m�,�xCv0�(�`G�$�'k�>�>�5�T��9a4�F�m�>*M�꒦k_��VY�t/֐�l�Y+S�}�!��>���x�U���p���:`"�C4�2Ҝ7;Y�t3&.��CnSƺ
�F̡0��1syF�o�uP�mѤ�}z}��[a�ДЧ�y���4�t�;ss�Ӝ#ņ,(aF�B�J�޼{�̭%Ie���&��=zB�|�?*���Ӿh�jcyO��Qk����n��S�W��6�4o����M* �$Đm}ws��m�j9Ë�z�[(<(�;`��x.{7Q��9�+��7:�ժ�0<U���cǗl��^���VV�V<~$�����<����N`40���fa�����(w#�0�Gy���X��
ܬ���ŉ����g�ݍ��>��Uf�G�hvq�do5�(�jo�g{/�����v��]ｿn��l��4�`f�+1�|Փ� ��6��+cs_��V{�|t�;�˱;�>�X���W�AVu�+�hA���SJIP]�!��@�H2��`����itQd��P0D�]�e�n�s��pvq����s��%ggt@f�t�8+a�FUu�һ⌍��*Z��^�\E7.�DϠiN	La�_M��ƀӹ�6�bǝ��I�^;��t�u�� I�-K�6��!���$]��]?��?��%%��M��-F��?uP�{�2��Z]�Fg����,� =�F�R$J�� t�@��݌�B�5�-5x�V�vF[E�,�P/Zn�����mugd����+���*�Rǯ~7F�!|w�h��=�@��5�2C���*��ԭ��]ZC3���ޥy!����,�!��ң�q�sba���-Ҿa�'���.sQģƫkL޵�gڑ�:},T�Y�kl@�]=�G4�DKt��;��� �P!�u��}�b�2�mO`��ۿ�fÕ��8����ӵ|���	��<�?�f�E��~K�=j��Xv[��"�0.Փlg�W5p�Ih��l���o?�UK�:�%�b����C
�/�/\��d!bv���v���NT;�zok_��M��eȟ����;9D���v�4Z��x,���V��L��H�����.
�M<:j�k�l���y��Yj�z��F�xnq+���������]�VX7cs�7B�+���q"�r�I$�'�]�WHм�ž��qt*�O~�?�����5�-O���Ǿ�cU�N���}���_�󚹅e����Ļ���ץw�%���v^0v�	����M;v�臿�	�I��=8>s�߈��� �1�P��?�U��$4�-Tj�3Ml-@�/K2`���B���CSϼLf�c�+;�Xى���Tdb��0�8��5YO{k����r�!�R��兾��b<o�Tyй:�?�r,7�t�F2 5�]�ddr4���V��y��!f����Ez��B�c4��J3���F��Y���KHG��r/���p'���\݌����3��Hi������9�v� Q�A5��N�	Œ��z�cq�~f�`7�T��t*�/v��5�7|�5����)�D��+;�$J��|OS��\��������_������e���$�g�`#j�?���[�����GWal;�@����C� �2S�e�<���;B�aW�ʖ#A���yB����@�ZY�'4v��c�+�]�P��Sp?F$����W��#�u~�b��;O�Kv�?�X9�и�rf@�|�9ѳ�g�7u8O���D��Bʾ̴��$,�)Rz��W)5dմ����L�������@2�W1������/q{�6����C7��;�����b��f�fB�4I�˰J�l�b4S��2iÙ�n��Yv���s�f�2wd� ���	�֙����ά�ӛXj���9q�}�<��qh���"��"yQ�����˳ �q~�8�w	��;�=��Z�Y��aGq\Ch�1�|���0��pv{Rc̢�HC���G�V9���(Q� ���u=_A�Βc���Ԁe�o�R��	�D�����еM*}�y�ݩ�\�O��m���=���MJC���},"O ^�v�$Po���"��	��B��O5���r3}NC=�o����r�x%�W@����E����(��%��G�=��d͉1y=XSO8���ob6�(�O����D�1����o"8Q#}oەn#J�f0�+Y�m���&ElUu��k��_o4����3_&�f:ȍ��)Ր���۠�qB(���<4}I��3�0�%�˹�er .�#�"n�u�P���?�Q4�eM(M�J<�����`,N�ABIN�v^+�&���\��&ZLk�]�(��>@�Dyl����v2^�O��\|]�.,kH��F��|�AF �і�y���љ����5=���$�A�`�'�3,I9E\?�C.<H]�Jl�0�'
y� �Z6*�
�\2M	�
vH�wъW���z�5w�oJ���՜��S�����	�(���dlA��f;A(:t=�eZ#�]��ޛ\�-�t�D]�Ul�b#iؕ���D�$s+N�R�kMik�(�)^�����%`:e���`Z�`Z���e�iN�0|�x63~Dچ(�/��$B��M
�qD��0��	l�5��%�V i���sc3��]_�y�[��!��%��r�F���v�/���Y�|�� *M���H��雾Y���-)�b�b�����0��s�e�=�TB Qu�D�����ۜ8L�����/��"Iw��+;QO�c
�敂���X���>�l�&8ۿ?�XU�V�y�:t�F's����y8f
��� ���Ѭ9�X3ª�~[�tP�Y[�g�鋃�)%^��ޢ�>��}�*P�JƏ�~�?88g�2����/iA r�h	9]8���u9�?��p=Y��#E��0/�͖KX�GU�T������LHq{�'��#k�?���kƢxD�Y���<� �Wރ9�goa�2/&�^N0����=Y�_�b��z���e�"���B��+1ߒ�6��n�	�Iiu����Zp0�痂�&�oZ����v�N���d�+Q@��#�MYvc�L*j�C|������`w>���n}X�ƚz�Z�?r���|�MD)mx]X���f�#��7n�5��K��v�-3U�w�����j	��e�i�����7��^{7)1|�4�(��o�gY^����:K\/���;YG`$C�HƖ��B�2-���?�-_�;n�DD�t�t����_y?r$V_�:Ҭt�w���������#��5�)c��v�5`_�I�2�1����+�T���r���If\�MJ�Od��R���-Bc��.;Ԋ$��a�dh$�Z���&�R,���r����p��,��6Ri�����_L��,.v����	��������fEz=�Ʃttb�fXW�Ku��֛��8�veH�T@���U5�d��$�YZ�\�f��v�Ch9�H\���߃����sD�>AĒI]S��PȊ���s3�D�#��#���x\%���h�GߧիA��	Q��)�paXA�J�kS�p��u 	�>��U�s<P�����&q�V�]}Y��ZZD�/�QaeyNh�j��)y����$�Ʋ�����@k,pL�b�p�
�Q?�<����+�:�]���m�0A�D�@`r��7X�ng�t�v� �|ȇ�V� �X�X�����=n�,7y����Q��j<�VC9pp{�T��}��0��e���r����f�'L���"��v,HP�oʺmNMV"}���(�"���&�K�w��j���_��~�3j#)�J\���?�O��Q�,В�L����n�<��Ȝ߀S�z�����3�?^�a��<2i�;G����L�ŔaDkWE�g��&'}pX��Zc�yQ�
 e����k�3k��j��x�s.�A�
�v�?�R��3>X�yB�u;���9�w��%�<]zC�����?y�h�4���"�#>��x�	��\m�$�&�&/x��+�P�]�5u%�p L�u�׎���M@g��{<V�x�q���<K��j����?2��M�|��ѿ�������	��,f��8��GX���zJ��Ȅ��$��h�ç*�6N�	�[@Z�f���e�0#3��My0�N�?��G@��f�̗}��Ͻ��22�aڕ5�Q΢?u�ѻ��"o'b;\��$YReZB��:zшac>�&	S�����s|�����`���O5��h��H�bL��8����U�q�&`���V�� �َlhy(f��e�(yq�{��$M�O��#������0��.l�NݢN<���c�Qя+|�:�f�˂U�	W��ۡ���hZM�Fgu�(��V_a�۴J-fӇt��=1���Ӓ�V�T\f"B-P�f*�o8�9�-uu�S}��-�vQ��C��:�ƕ�1e �u����Q�o���sƉi����C���4��d'�Q�_fM��x-�<�q��kd��'!@�F3$��oūR���4;���B�_����R�������VK���귏@�a3�!�\y�b;�}���LGQ� �A�����Y�B2�G���g�C���H&F>Ib�t��vh�9��(\��2o�׀L`xs׵�G�w��.��} ��=�����~��×��tg�U�r�b��m�3DJuW�%#l�NM��u)��!��1-���L��C
��ex+:XB� �Vi��9W*�n��G+֙*���J�ɒץ�l��,��ǘ�Y��D�Z%���#����������>��H�T�7�F� \"��-�%�&��.��|����vT``���`���Q���ċ2�Ʒ��;�i�)���=�#�A9jx����s@4��^YI�b�e�"��C�����'`�;���H!_F��w�01>�<�t}j��*i���o�7ܿ��Br���05ir��\��oq=��\��V
�-����f7�GP���0���Y��t��}f۫ڡƏ0�g�Vt�ò�P �V����,vK�lf�˶�Y�,n�Ip�/d�*�?�g� 
�M$K%�*s����oa�\�;�g���'b�`���/���W���X?��C��\ ["��Ovo
���5IH�F� ��k5���q9X�p$��u�ҳp�U�#�aÊl�Q#IQ�V��l�#u�fKw�S,bPa���ZU�A���R�B,Q����F����Y$O�hB��kI�d��ݿ.1�<�h��dE�yl��7d�'�e$uo��/�,J�KȀ�A�zq�B��uP�pa.��(�u�qc9�n��.�{4��b��}���g��@�ѯZ�~��5\0/���ޠx�*�f�����?� ���X�e�ĭ"ԥ�]��T��$AC���дLH�U����;c1�:�����mJ��$V�D>�������
/��"S[��#��Vd�Ī�#���9�>	��,�l�v]����*8Z�TD���b��:9��S��r�n��w5�S��ɜ��m]�dR����5�%`�!G���N�w�6h1�=\���,^R�UM�����U�Jٴ�g�ZK]�+��D$�m� x�����6c�6���3'B?�hM;L��!E�ԯBBG�$3y�����NЏ��3�����;{��1�t��Wl��hk�4_�xB}_�8NT��(#��G-�'�n�	��m7�� ��5Qa�y����������	Z܄�p����B?$cNά/2���Fgs�U��;j�f�������t��y���8)�+�2���&���!Lm��T�]��?i����A��B�]e�'̌s�J3ȮS/cr�ՊB��!I��(�)������z-6`p{�h�x����$�ב��J��&�܎Ѓ`�n��r�{=����{��2|�]��G5�l
�%���R�񚷔3�^A���3W�<Y3���
ϲ���e5'�f��'�%�!�COKi���|G����mLRՄx��R��'��L�ͺ���/cy�QD<�#��[J�X�M� k���3� �EJ��c�q�4���:��^�����?7)�r��h߀�U�?�<,�]��*`U�B-� ȓ��o�M�W���2-���*�Hbc��:������"o�F��n|IBN"�1 Umؽ�x�}��aT2�6�vϘ�Q�w�5��!@c�UQx�X�R��5��"�9k�i�T��GBpm��E`�'�;L�#�(4?����0�]�.�\F��B�8�+�Y�����GxI�$�c������C^�r�!�"��hh�Yz7E�&K薚ѿ��p�$OI)�c�9��K�o�*�{å���ī�p�^�Y�� �>���A;��`�zagF*�/2�l��w�t��^J�EՆ/��au#����ɊFF�n�5�1�����޸����� �C�d�N>����kp����a|�00&���ŏBNO�t�h�j�Y&f�K�z����h�2�礻1w:�+�ٷ�ZP�맯SH;$���	AI��>r���B*@ `�f�N�$��y�����eH�)�)����2���lG%��mn �D�T��K`(���^n�Z!������ID_�o��Ϋ+�6��h$:fT^��F����>�--�E�B�G�f��nC2�2�&<W��6�+?��{^7�Y5r"��+!銭;��(�q
B^S�Nì
S��F�ڮ~��GK;�r���8�ø�,�T��%;�s=6<9��X�xf\F�+*)7Ҏ��q�Dj�?V}�_�RW��# ڵ�fF�?=O�i�L���ַ� �����d�h}�3��!��i���K����T�a1�:c-��#8�soLE"Ef!J�A�&No�{s�@�fa��V&��(HX�³p�݊>�1}S��ZJo߯����b"c����\8{^f�"�l���xp����!_p������1���N��Cb�!%���<Fo�&(%˔�Gs��}O2�����a��$CC����b|��߿Ov��p���=���`A�F�u,lF2�8�������!�&�g�ֆ�a�C�v,�.w4G�����\f�b���3_���@��ݴ�8�:]U'GqFMbd��X�e� �\����eU/$������IyZ�ظ�l^�+>���Hut��©�]���3mxd~����-1f�;�ݙ��ƕ���}!t�tD�m7vC����%|@��г�3����w���'��KY�.���wI�����DK��F��Y�_q���0�Qp;�r��%�6�( ��ĂN�(��J1�p� ۜqj�8y��QE�Q
J}�pn��J�|.9#���S�y\�G1ݰ~>��h|�ފ��zy
G��R�=G���pf^T�.��3aT4�A
�e1 9W���U,��j+	׹�\/�$ըߜ����VB�q �"�5�M��?��Z��U)�{���a%U�aCx�sj�i%I�JY�kB�Ɓ<�����ֿ@=��)��|�)��	�U��]®�.|Q}�1[F*o8���l�g�SZX��&\{�D_|���x��KR��;��)Eh����}e^T����A2耡��i��e&mq��O�w��k� ����k���6S$'E������)�E2��|�#��O!%��V�A=�\1���9JV��חn6��T2|�z�`yu#�
�2���:H�Nj�U�������
���R�i8�[�1�&�?��ۯ�ƝF������8Zju���@�~��У���������9�S���M"�8z� � N({j�8h�3�B ;�����tj�>I�=���{���]�/��ѷ�6��ۂ{�Y*�Σ���)*��ě�劄�
�3���z�C�G@ᣮX��Q'/�O�^[��"�a�9�5Y(6lݟ��|���B�B�k;��6��ϊA�g�Tg=�+�3�����q���:���{˳���4{�Qy��l��S��Ա`9�����/#�EJ�)m���*$����y/˵\��+ʲ#��C)�>�j��#e����� YXs�p* �vK��ҕ�R�|l+Q�I?��5��D����`Z��4�|m�aP��\i<	k��A0�s�K��������7��R�t��5'ǎ�`��0ҶX��,��*������V��T;~_]�@�m!�D6�Ǿ�{>���~1e��*,/5�����'��͏Vu ϼ��o;���P��~䚶�	Wy�����2���l��k��*p�n��p������q�=�}-��=�����~f�8�Vƽ �x���s�Rt�b'$m�;5��|3)���"��Q.w�ڮ_�M�mֶ9�|��|=8����p���(��˵&��{�=�߽�T�:ڎXv�F_�p2Mن���E�!�P�G�+�^�qh��md�^:I:���N�o����4��e$�?2D������U�E���������x���mɿ2P��/#஖輍��p6�Č^?.t*����|i����"�)���_Hߏ8}��f5��@�-�F��t�mčQ�����>�@�����'[�� ��]����Xy7%u�i�R�&��'�N�ÓA�2�1Au������7X5��q8eH�|yڢ�Ʒ
�q��s>�&�vٝ�Aը�Z�ss��Y��aզ�D�L�;7QP"�e���%d���jU��]� �
ˉ:[ 1��-|^�o�&R��9Z�u����G�������^k�o9���"�R�|�( &!P��	̃��*��j��ǽ&���ӚO�<h�,$1���� )u|��Z�?�GE���҂Õ���45o�4(r�6�a��.pS�{'o������[f��aDٞ�;�a��Ā���n� ��J��z�5���c\c��&����5�U�2��؍��c��A�����Q����������Ir
*�vg�}J.S}��<�,)�ض.�~���=>ݫ�(�����Ƶ���=ߑ���̨zp��%Kt��R�>�ʢ_�.)��NZD�C�����>���B����W���S�y��|��V�<�0fl+�u�
	���"�pr�	�i��!3=տ�Fۿx�Lﰠf��bB���@RT�ʱ�ϳU�;z�T%v|���e����;�9l~��^��X�����&��I��Yc��|��̄�}7�eT^1c�I`�Yv	
���ê�:a���ԛ	����[_��Aj�R�8��P������*N%�m����3{S,&�$��X��w���'�O�zu��3��(���2��W��ǳ[�SL�)[V�
%�M�	���^���Nm��n�7�����	k%?�<��>b�4խ�����g⿣���.ie����U;�)ނ@~@�uk�������Ozs��ou��*UD��c�\j��^+�����Z��qW�2�+6�޶��,2��ŷ�m��sa<�����8J
q�\d�2#�sB����9��9��"u���qr���S�s]��!z;	�D�bY���HK^�p'���{��q��;�qc�xk�%  �V�T޴x$���⻅V�d��A�
�z9~n�9}r�4�0���^�ɽFX���R�S?
����O�M�`IĚo��-���'���������'[�v���k�	�l�}���^�I�xMOB�PE0��6��-"/&s4A@D�n�����dע�N$l;�G4iI��	2�z�_�}��u����/��=�BHD ��!�x�x7�1���A'-~P���Hٻ���n��@3{��6��'�Zz�XH��Y��{/Q\e+ �7��Ŵ��.H/ܷ.�`�:$)�M��is>?q��7*�����W�.�@��(�7����~u�)�i;[��vl|��Z�!S��?�Y@�-zT2��fwNL1�ü��R��V+3��qJ�����0��!�S������PY�����?�F�Z�"��Q0�x+���o��~���`;]��W�#{ޖ��>�6�=����U���y6`�W�p=;7��k��#���[�+�F�v^p'�u4�E���m'=�n�1�0�G�����Я-��ǣ��h��d�r�Vґ=�������P���S,���#���Ͻs��2;�Z7�J`�iԳ���A�������r��}fa������aT0�ܐ�+3� i�h�ic1��lO	��H~�&�h�_`(qm5�C�7���%�:C�8�����"�Ȗ
]ǳS2�m��"������rO��6U�J`��F}4��K�E@~m~xE�"�Ra�N6eS�,�%��Q���;�{�U��a6��� �J�$�<-�I�̾]N[�ؚ8�\�J�vlv^V�V��pEl����.Y���]���nL�����P&�v���掞-��KR�Y>I�eN��G����P� ^�o���^U�*�8�\�K�g���,V��M�`��r�-갤$������z}�T���c;��I�.2?z]���l� ���	��+x?���Wj��)��)����jP�.g�F��lQ��뇢�5�	�J��F]��V�*k@�}�<X oW��ҟ�������������cP���cO���~�.��a����@}�0�>���C���D��>��	u����
H�
d�`f���$V4��X�Ac�~3)��iT��I��jrO���N1M�5�o�M< ~r�&�x�L����]�*S��'�sN�^�s+q]l/v��p ����y�3:.��S%a�C�[���%vK}^Cf�	�� � ���	�*n�Ǔ�vؚ8�i�Ja܅D>dR�r���,)�+R�ƕ��i���k�$�)�瘍+�Ģ��MV��"���70�-�Ʊ��C��r�{���kU4bj����>�5D�[��̜���t)����Q=+���(���|T�+�����m���Mf��~I�a9�R*�^a���W������`��vk����v̋�S���;j|�nGS�ԒO��3E��Wt�ي�2�@�,��ϟ��K>��z��x>)T+��r&&�n:�H� a����&��s�����BN��e���j �iS�cܜ�����R�2"y���ɮ�-��;u�:���T�����k-%O~Ld�-f�W�K�$Zx)@@��䣚��W#����B��ɋ���I��Xfq��U��Y��.ս�O����'�M:�C����Wc��7
H?/��"� ގ���}D\��c��1�����Nt���2$W�Pa��3(v6ix�5���KjN�P⾚���/�ʋp��W��zw�E��Gv :���D�izy���j©���/h�0�d�����Ea�&8p�H���3�{ ����+|��>��K�BJ�-���ǭ䖏0�U
i��8nD�{�9M�CV-�Å
��V69-&x�E��Ǘ�55K��mOg��K5�a4�_�yT�#eT�S3�@�ȕ���g8��俪uSMe���A̱��=p�h�G�L�+���f�<CA1�]<}�i��uon�e�M�������dŧz�����D�zze<����U�p}=9�Z�]�t�fnWx�+�?{!��!���h����S�o�_^`���uO��\u�����X���߅'$wO=���x�4wK��&L�iFن��s����˚��
!k/���*�S-���R�P��~|K�q��Ž�ۊQ��>SHH��]�p�Uz@"�h3Eŏ�����º�`�D'�7�@����6������,e�.<�����ǼF�NO��j��W�*Ɖ����K�G�H~#L��HQ��*�	�S��m��lL^�kK#!J��C�~��m�2�"!����ʱ s4�F��t��ݒ��c�I��7����'vu)�c�H��U��tv�('T=��&�f�
.?X9����?�Do�%!�Ȫ��S0�*��F�)�����6��7��8_�-C ���p��6E��T�/|5 {i�`{=_�e�E��:��&�B:��}9��a!Z�@���_��"'���E�?�YGS�������e7�﷣1-jW	n���t�4��=��3�Ǽ_��٥�g�����4��R�%ظ����*W���=�8��a��ĝ�0`��Ć���֭���.Np�+����AW�������_�i�*(�t�H�=�z�K�I���s��@�I�K���ї*��cЂU�(_n�4�*�J�3G6�qGfm��Mi�l��xt�R�\0�]u7�#��Պ�O�. tf�ns�e�p���hJ��a����neY�݌ҳ	5�VA�	����������ψ��i�ш2;J"�5���I�<f���DI˫i��͋�E�/r��A���E7�B��<�GH��T5p�fn����P�!~�<43E�ΰ<�[7mm�G!l��ÓE�w6����pB�4��8b�H�ǆ$|į��]�>�Y)���_c;\�M��fNm�26�:mW��7G#�pY�����|��k(r��:�'�J��5�u��%��/	��4� ��~�GB�`��%�z{�My��l�)Fkf��^K�Ug"2}��0i�?���s�7ӊn�_Q�*��$| WS�ex��y�p��q��
�O�P+m$�s��@T<��G'Y������o�fgɦB$!I]�9�$4���Cܞ�6@R?{m?�[�)fe���{ae�hO���5�p��-��yx��\^?�����K�f����Zx��i_�e�ZE5��I�g��D�弴�z<\���}�wP����V�����+9��G�^���4"ƙ�T�*�0ƨW��gG!5i(#�l�5��FX�.��-!x �v{D��%r�_^�ӊ:+��̺u���i���r�����U�i�������h8%{l��6|�j2�;&��s�tt�+�]�yl�_'$�>�m<�颿�Z_������G��~���2Yy&謷�!�ղl�n��t�6(�j��7)��g��}�F}��mi�C^d��ꨴ�Ξ�E��Z���_M����M�/�W[we1?���i!}��g|���S�A��Y����Z�dLF��{k�,���e��mޫ����!s�Y��;
@��Vzs>DH}��]9�Q	kQ�fՙլ�y�vG)d�.���^v~�B	�*��S�2ע�wm<�[�9D�XU#�^��7&��]��qA�vl�ғ���N�[WW�x�-��i*�Yw�\�#��;��K`80 A��\�r����*���`d��d�V�I�5�cQ����<<�%�K�4@�]�f� AI��x�o߰gD�N�������n���i1,��f��nIZ�1������9t��,?vOfq�����2 ���:�Q���X�S�W)��~.�t��2)S�}���}l�W���z�7�J�BY���_@�	s���nV҇�}��Õd��)R��4�]ɾ)�(�Y��p1�zk�B_r�KӀ�6����<�����A��l���O����� }��b�w�WDF��I��%W�}?�9��m����N����Z��Qj's���Q������ęh�LH/�s�0c�+�!�� �́���pXX��D����~�$bg�l�0�� �4]��m�������K[�^�*��v2$�鷽l��P�4Yp��V��ZQP����f��iD��c+��%K/J�@�M��/ݴ���t���"T��E�`��L���k;�	Y�t8˰:L�i��j���"��l`�Z�լ]q,"0Y���nq�/rFI��<���6/T\��:!�mp�֕���^�G�ժT�>���ٯ눳DB����}�i��e)��C����\�_I ً;7B�5�)us���(ja\i�P>U���(ś�Om�I�x����
���	�%�G�+��E�`����P�7�Yc������%�nh�O)j�m��y/� �뽘�S�u
N>�����3��H��#cMxx�*9.��������p[q���r.{~��mZ��P���*���*���_��k>�E����=�U�\!�`�^G � �h�@3_J=����z�����4,�z��#���f�R����b�A~Qp�i�V~��=W�f���i�:?(?�`oߔ��qww�l�/��. W���fk���ņ9�J�|>�L��E�B32d�!���*>��#�=�V�"3��T�O)���%�j�㵺'X����(Xņ�8s�$X"zpκ����B�E���M!jL��z�[|�3��z� !>4bm��	`��n'�W[��]*��$0����'�(��,��T���?���X���YO�A"�_̸��z/����C��8��hm�A���PN���X��	�E��;�
1��]�3�Kn���|����8�5�fj��}tP�gI�'����`�}Q�����m�y� �'JLN-�o���/f�;�'e�*�a��RoOA�+=��Q�nGI>��?Dg�=���` <���25
k�t��1X��ɿ}�c���ţ�>�������/vz`�C>���^r�n
�p�zK�O���ZS�2&��^�k��q�����N/r�jSG��ۀձ�w*��5.ʬ���7#���2K,����>xvuc�@V2u_>f�-��g[1
�xϦ+'��9���l/�ØߣTI�-W��6a�i7<rA\tb�t�Gp��@g��ә[)\�`��ۀ�N��3U�״�)0�W�[5<׿F��"M��V��u;X�N����&�o/�
N��D����)֣��:HUᛖ|�����tZ�6�Ђ,|��;ш�|{֌���J���1[�уS��.��"�!�����@�i@	�}� �v� �Ǫ�z�8��~���[X�#B	V½CC1̽�}��ߚ|]rC���ڧC�i�`:�3ff1$�e��T�ѻ���o����v0f���h{F��8[`.�/�V���~Q��}������4o�c��jWv�^�pj��S��Y+��O�]^՝�����2��C��Q�U[�����&�>��ز[eź3�ߜ@_=䵊����;|���>p1�
�r/��X� �|�j�!��Q���r�V��?�(����Ae���ۤ����ǝU�śȧ�t}2����_�CȻw�BI'1͐���z��闯��	β�ح-{3��v6���W��ݤ�0kmG|R��w�M-m[h�{�=����X�)VV�}�H�9:z���=d���⾺f�df��qڞ�L������m�.v3��(�O�x��Mg#�h��}��SyԢ�Y�0���w�,<��Cǫ�ZU)����GK�]����+&9���i�8�^(���Y���5BѽJ�:2��3j�l��<rW2Er�'��� �a�:}lp���͛���B^⌃.�>��|l��9����p���Yd��O���qik�j�=^�6WT`x�7����{��<�]��x�1u�6�Q��v����� ���HQ�`:3K�҆���LDpX��8Bܢ]�w�w3E� �_W���X0yx
`ǹ��m�x�e��S-�Lo�^2�WF�H;0 �nwUMUs�e�p ��72���,�T	��IE���[Ӣ���_�$�p6Y����G�Y12m�@P�=������~��f`�f�anw�����j�2�/x~=�$�k��(�����Ը�r���2r��f�SIc�:�v�������v�BR��?Fq�=���IT;�h�''Ԁ�Q�
-8T}�sJ�8�ϛ�]3(2��+�E���V�ty�4F��Jl3<g.#�h�ԕ���C_�>4�%D��pf�$�y��ծ�������c��\ۉ�sg��m��q��J����o����V/��Z�����
�u��>�����y>�C^ўŬIO'��4
�g3u~�]���ɖ�_m�I�;�(�
�,ĄP���[���8$��/�@�%��x���E�u�����J����Ӈ��;�� �BjN��8��h�%d�	Ǣ��\���y&�:(u�'j��ds.�M
� �ܚ+���Ð+ǧ1�q?��Rc��-�Sv�_�Z�I�l]�Ka���o�	�����؝�S���L�kd���7��נ����� �'/�S�Pq�*�?��YTB�Ms�ۚ��L ��$�2�s�+V�����&_���s�� ����u�M0cC\k�u{�����\�.�����X3b|"�F���szHW�Ӽ�pQeq�t^4.��.�'��)�������ɡ���gX��Wz���۬�����<"��{���.��_Y����HN�f�{��Q�=�p��ÐV ��㻜�����x{��=|�ж�����4A��^c&�zp}J�?��o=5�'h���2$��'F����޹������-�!����i��w6D
���I?�,X��ȁ�QUs��`g��{��Y/WGŵg6Q�Fg���Tmeu�y�� ���Q���v1�[9&��e�/ȳ"��Kn�C��"k�?�O�����\���J�p5�OH�yQ�Z�0���u:�3�Q�]q�Qd� ���;G�v�^��RO�/�zˀ}D'pL����>�v���ļZ��(v�L)�����]��῍����r�4*�_�!\�V%��z`ی���|��Oj p(#'p��{hK��n�,�>� ���0��G�u��a��g9�_���y*����*�n?��I��u�l�Z��h�����Q*��o�!�}�o��3�j���	Ӂ6�"MCl�T�� \j��%?���V���#�`,#��j�fx �uo����j�2�hu�����d���!�&�j\�dO�8̎�����F�m�?q��|� ���7�\���D�CI����[#N{Wh���S�egN���tI`c:�U�A�E�k��T~�Y!}r�w�Zk� ��w�0��ekRa��$��ZD1��ZZTT�C���B�kԋ�I�n ���|�8[D\��1�^���}�G�}�3�(��l��~�QXb��ԫ��b��8n~�O��ã\y��ӿZJwT/Pb>��=�a�G:!�W����U���E�Ú+r�:���?�uV���i%(��P��guٍ�{�9f~-	�jn+S Ѻ�E�%J{�TU�oS�>WQ;�ĕ(ڻg r-�/\���R��WSY�@-Qܔ%+e߼�J}y�%:�Z<[�4<U��ئ������>q���2K��R�6�B�S?VO�q��|������йڝ�K���;�>!���O�`�='��ԬlZ[M"ת�������s+~Q�ؾ	~�~��	.M���|�B�ϙtt.6F�:�l�#�.�(`�_�K��f�,���G]&K�]����f�����\j��_�e��Qg�ww��S�q�.KU^����I�^w�?%.C�5��\yGJ7��� �����P�!���%�NQ�#�ӫJ�F������V�[N�^^�:�,�uF��˕G�>}�P�/Y��ݜ����QmW�;GFH`�BOk@Ĝ�
2&��ʊ1	l��S�� -'�Mވi�2	Eg�o��y@ș�s��Z=M�Kt�'�(���l��r�u%������=��(-� �Af[(DZp������'�R+|B9�z�?L�kף��p�|ԣ\�#�K�F�~�\���1�>��d���=������l1E�l���kd�y�X�d�2/�c_���p��[|œp^�v�*h=g&����̻�n�<�����N���T�/�x�
�u�!���ZH>���d��I��ߡ�����-�H�};��|p/ K$�Ы��Fƿ\M��Ff��\Ю�':�rSr���H����<��2�S71�W*��=��8�v�a-�S(���2��DpN�^ސ�|���&�'Fkd�2�ϏR��2.Kg���%�� ��J[��b�2U[�Vv�������N@���uh�ԇG=��D��wkIW�x�[�ʢf ��tq<�S�'SP�����4ֲ�#ɘ�$�fi�s�+���3Ǧ6����6�-H�V8J�_������:J����eI��o�ïtR?;LU;c�.��?�kp����]�V0�f)®hh��U�]��$���fy�����k��zhs�1E�@�Oh�t:N�d�b�>���ȵ���-9ȫ2�8IE��j��(
�vh�dTQu���Z��(�OB7F`%2*���0�Q=_�RwJ�{3�� ��\����ɲH)������Q� �����V��BI� ;�x��(�@#��'�U1`������!�{��Y���S��,�M��9�����G:�D�7�q�!�F;^�HI�����~0hZ�l��T���<j
���ؠ;�k��P(B ��#U�$���gc#��UI��	�@��x��T�%n	�M^Aj��6��a�|l��] �C�g#0�?b�W�����Mf� ఠ��K}a��^�g)�ܦ
� ;�q9���'[�Ɉ���*����l�%lo�ͧUBf�X�f�[*�N� ��u3�uS� ��X�C��^�3�x?g�	_�e�����/���G���CQ/�<�R��Vi�KS,��wзB�x=(���a����달�!��d��&V���Ha~o�ʟ@:�:^��f1�#�s߽����'����i��o'��ZZ%3i���M�W�qK��D������q����@��*����:c�d忇鈿q�ش�	�(:�7zF�����.z�m^�y�r[�Gj@�o��XlĠ��_�pU\� uD(9j�E��	֓��;'�k����?6����V%�4�9�� �L��`=;�	[��Q�S���$����nhcT��/#l%�Fs bs�7ʇQq�� 5�/���(��Z�+i�m�����F@�*uk�=�j�zQ�l�YI�ދ�o���%�_�	?���`��/)S�S�8�\�|��lجS�h�CEbk7���Md_�����,�>F�_Z�
jo-�̝^�L^M�;�t��)0�}u@��Hp�y�@�DeS8Z��w�K�2����m�~!����cXw��N�*c�[UX�U��� N4H�Y�ϓ�B���2��$��j�$���'*��d��j���Ʋ��=�*�5�9ATK�Մ}�v1�_����s`Dg�$ס�84�yk�/�H������d��5V!�x�)�kt�J�Ymqτ�*(�M�!�em�V�����@�	� O	DFQ�Kf�^�v�$!����z^ۻ��k\k����J���;*GѾ>���PM���?ҿ��M_N �6������B�Lv�ź�o�9�iw��-���<���~T���IAS�n7�>C���qF�utGo�����3 H��F*w$D�����2�y����@Lo���"�%M|�,I}�h���#�n�;Jt�+�W�b$K������Ĭ��BH`��hd.h����L�Y'_�Äc��:�p�u_���oN�Z�>��;I_R�O�y���:u��[|��n�~٪����YeQ��|b��Z��l�)��3bDt*s_(cg��	7x�i`;��k2H�_�n�]o�JmD�Gخ�Ab9S
��"Y�xhȵ��T"����������x'�M�HC�δ-�,�4Nk,l��n8�}cTC�o��pR��h.�,��(��B���6��?��X��nDR��q3��X����2}�rz�ܢ�Ԭ�BA�K���(=�����P�(��I`�e�V�$Zj�r�$����3N4������aV�w�ECv��A;ϓ>
�@:�Z��<�n��@�۞��h���Q� ��pnG?��Q�(�)��d4��n���Qwy�ȥ'4�zJ����Ԕ�&��&�7r��S&�T�-����T*R\`TS3y�i��:�B������Ԇ��R�`�ڍ���+�ew���d�L%q���ת>5X3�6�T�CM��s�moYq�nI9�đo�_^�X���=�g4ե���|tc}N�Iܴ�r����0�+`��'R��c}����ԙbM5�Q霚E�CҊM@��*�^��y�R}9���F�U�,�8�z^Mc�~��@��~�lSϻp���!F�ǧ�)V�X<M������$;����4&�8�8�{7]�t��
��B{��9Y��2p�@����FӲY$}ݡ���<��<L�OMk��M���SW�?�k9"����h����2�w'S�Α�uau�u�J�Dv_Ը���d:��骅|�MA+�%�Jw��.����E�
��kD��%��� ���c M�UfQ
ձ�5H�*�N$���gh����%�f�0�����&�@\� \�#����ʧ�,n v��"�u�jc;u�s�T�"!�vn��]���>q��.zy���Ng���H�%`��'����J$���G� ��J�/
/���w]�/�@f��N�ic��w7��(4�$	�&c��Y3�W]�{ۊ�k1}�s��ɠ!���iF��9ڕ��e�4J��(xx�%��P��Y�P��Ʃ��0��v��#���߀���r'�����ɾ���F����'� �@$,�W��&�
���g��l�T����G�&��Ϛv������R�yX��gDB�ES��z��e�wM^m�d���+�gÔ5�O(;�.�UYn�Z�K�r')�v=��ɾCp�B�z���xo��'�)c���W�j�!��,�ҍ���˚�;܅)�O��pW�ƋEv�Iv���@���!7G4�'�=kNt�V�e�˰��������A8�9h8���3�`f	�#�����-RRT�Hi��q�ۄ��*:�.Y'���Q�+�ט1
h���5�֘�vǜ}e༼r�1A�7�N�ݣ?�%T �;��������σ�aa��ֲ0���|U�o0Bfc�yFF(xK�����{����ӏy���������d�6824=�C���EAt�B��y�jm)��ѮPI#o����\D��H�,�i��G4ɹp������0ف[1�W&a4J��������G�'���G�F�o��2)�pl\��E+؎(�h�ě�ӝe�2���pRJ�'����n�;
�[����'�'O�C�T:4ߘ�׾jzrV�*�erb��g�-�ډ���^�b�S�4t0hb7�� ���>W?��	c�a�D�/�H����F���E��{�,��άz���ĳ������ϱ^�@�K�+]�+"�0	E�2Z�X�)��*M�imn����kLܾߡ�3Bt-�%^�ښh��������ov�+�>h�e�/' ܨ�������T���D��ʞY���������ԬP���#����a�e
�/���f��=|��I�9/M���܇?K^�-|�+�In����X�m�?�%�3xӳ��s�W{K� #�o-1m�q���t�ur9��pf�b�/³P1�Z��z���l�GQx��m�0ʪ;��HO�4��;&��u'�$�"	��L^j5�5R?GM��(���4AS~�jb���{0��@+�� 5�\)�蒈 �,�϶�}�-H4�\��^����r��~�"��J{��l�nT�)�\�(������ϲ��Qf+8����_H�$��5W��z� S�3@I�IҞDL��:`CU�]�p<[��i��]p�g/�ٱg�ݏ5�H����;����Զ��B$��̯�)����U2n -DN��~�ys�&�����0��-��1��ApV��m�:O|i���� S�x��cy����u���/+�*�:)��Z+�<$�lǏ�C�_}�u�ImU8 �k�u�{4��P� 8¸�-���}��Ee��8�<e,[�f�*A�(�E�r�%!F���/�L$~�Vq�&Xj�4��Z۷5�K{;o�N��(�U�����C}
={��}��kWq3.�����>��2��>_ɱ�a_N�ϡtGW�Nư$�������U����$O�7ߌ[)A;�������,�0U@ ��r4�rP
{�>��p��v�����%��b��������)�=����F��)�n���?"���aE�@��G,�*+�e��gu�3c�H�F|�LgQ$���-��'����E`t��W�X��Ქ���l����%L/�-���ߍ��'O����MN"�g0���ր��E�w"S�B�D��]�'݆]qޟdK���G�|�	GZ�s��L:�St �+���_�L�c�ћ�1��(�H�-���͞cp�4�[ma|��PlO��~jD�W�b�+('�^�4�a6N&h���;(_�S`�O�tt0�Ա��u����]W�p���u&��{��Y!j�{:����S�ێ|�	���W\��Ǟ�����pe��Ύ�8��&ɹDu_��j�j1��T��Ц*��	���+;��m��M̸֜j�7EX�ȫڄ��T,	CRq�)Z�)Y	��Q(?��^�βu���W,8
�H,UU����橴���Ѻg����倉]"L�1M<��z~�!�J'��|��U���zC��1�}��z�&�����J>6HHO"�h�TwD�Z�U�m)���0tR��N;��Si�}��(��`���aJ�Q�=�#{�{Uov�<Y��LI�V���E��YT��	���1���xb}g�0���I�:�m��&�6'l��_�Q+�)W�-c�`W�xf[Ec�5Y	_��*)������l8Nw�P�J�,��N���w����+^�G���\t�"D��R^�1���g���y"Ex}Y������e�5�g�0�}v�%��?�.qM�9��;��w�H��f^�H�Z���c O�6+L�int��t��2`d�?} ���HYԬ�g����Wrh��r�sX��&�	~έE>E�\I"G�J��CB�fQ5
�k�k3w�}����"��6>z;�eT���2|"�^�Q�����@zCJ��<#�ې�ax���A,`�N��ܛi9�A����Ҥ�:v�hB�ך����Q��5Md��i�L�/�Vw�� R�*��a�p��b����.5�ˌmN�|���
(}��>^��V�������ۍa��gp@v�c�I�G�FAzL��j�ߔ�'�-B@{o��c��v'X����JW^��@�:ȗ�=Q2�SN�ɇY� =��G�����N�հM
�|lD��ӈ���̔�N΃{k������|Ǻ�+�A���,�Z���25�C	��]�=	��'�y�U�zz�ջjsB�/^A����6���Rm>����z���D9>QA���"���erɩHǮ\HeB��l�z����5��9�����
&��)$��&���e<]	Q�}���2%i����la��D3�`Vu=t�ݿ#����hw�M �S�vFVN%�V�d-���.Pp����cZIXl��-w��7S�&���)
N�ʗ������	��`���n�>i�~���[q�TB9����*gHkm�ݛo���a'c�%Hv���g�$r4��uDw}�_�C%U;�6wՙ�M2oAk���vn@Z���ZpV��F�����Uɥ��z�fIdR(��㡹Q�8�����P�?�)��@<���w.�}�^L�W��]K/�3/>@��hZ=�{9o��pҙ��L�C&�c�b�0�c�C��h�i�Ƽ#�t���G@*41��m��:g"ĶJ lYx�pJ��
�P��e0���m�'�	�������Y�5�QP��rEݲ�j���Y�?B4?���F��Ń�yX��v��dy��_��R�'X�?�F���Wአj[=�`������.Uu��;He����,)"����Nu�>O��[�g��	j��߹�}���)AE8��م"���n�>���e�*�YE�#�o�5�Z�qd�cV"w���&�~u��KM��}�x����J�CVK<F7xs�׸R�+i�������^#������2G�]��ۻ]�ps �)�=�|�_�K�e�\[�Q��2���q5ܧ�%��CQ+���V�K}����m�UU+b�[=�C���
���`Б[]��<D�C4]�����/�����q�?��q�:�-�;NI��IfX�s.�I\��r$g>Ù��n���Ln<�[i�6���m���>V���0���N8��D{�/~qG���8���rB5��W��Y`\sy[�蟡ˣ�)F@44=�ջ��+h+���K�y'l�*F$班����U��ѝ:"�&�i{%*4>���L:O�ԋ<��T ����K��s6 �7h��~�pk��t�Q��Ũc9q���qJ�0�L乄o��\$�D�Y�T��u���!�����4��D����T�hS*e_�]BPp�Pew�5����o3-ff��5�W�]~�(��ؠ=T�S�q!����z���^�א��ϡ�twH�}�n���K&4�壷����j��i���]J8ͥ��;��?���:v��}�.��8|�뼘3��Y��y��=��p]�I1K�}6fT\���9֤��fp�rYP�C�P��6��kmh^���ůg.�XbſX��V�{���e37�!�c�⡿������R�ɕf�"[��M�3GA�榼��ϟ�w~F���ۜ <Sk�q;t��F�r��>$`�Li�X���cZ�˧:,�	��R��^�ف.J-�0z��b"7n�SNr.r&:��|Lq+&�M*+�^mDlG�������B�����#�d�8������DpӑM8����S-�hq��] $+�Y��x�:{.������f~�3n�;��-��{��P�w�ូ�\������)9EƘ^u�)({C��,��<�ض�ިe�^=n�:iW����� �j��J]�r@011z�o���$��V��+��4r�P��"���M�d�"c���|U7UQq�ww��������A�N�{[�W�¨<�*ߴ���f�w�N֏H�o�7����Xq4��ai�v��pO���b����IׅXḿ+=[�n6�V榗�nc�����[a�����R�e�]������1��9����t>c��9Q���_IM/�M�N��6\-Xj����P�ulxB��%$��=Tt���a�h�~k��a5�	L�fs�%c%DMxs�|Ʊ���pؾ�{�F�) �'��,xGŸy�ׁ�,'oÏ����-	�PN�#���v5��}��Ss�i6F�y��;��8�^��8�p+��$@+-� a��Gx���"�D��nԱo`�A�@k'���ވ{���7�jk^ސj_��Γ��#�8�0P�@<W��u%�৳�j5�ң~����w ����Pb��]���@�*ߦq.��+�G�Q2�>�f^� Me��f��1�88�'���ˍC��Ph/���b�C�+�'�7�Bv���bE���$���h��j��R��3v���I�E$�6a�+ /�8� &q��{>#�u��,8m�U����q���Y-��o��8�B��w��B>ju �ӳ9�TwF��K���05oE/�z�ا3g*#�����l����8�SC����e�7�sa�P�|�/r�������R&Ƕf?.�[u�ܐ��dc�%�n��
��|�ࢾ"�������NSI:���o�7	]l*�Q�:
�wnssV���+��<��/pv��g�+
*,�����;����)���Ÿ�5NZ�$��T����mp���=��,Uu)iHe�<����c��Um\�8��������yy������s��7v�e��f�+>4��P�7��h�D��lh1����������,�����{0�upe�o&���w��ne唸g����}�F�S~0EUp+��,[~�@�J����\���*�K�E��@�mN�O�0���0(��!}�ߺ�B1)���C�k0kJ)�S�HDÄ]ݻA;��wq�zJ�Q,�݁�2�T�C��:��D��)&�������*�^� �QG��e���q�Ǥ�+�O[Tǈ����F���ڀH>���a,vO��ZiCa�@�<�r���	��Y`��Kf�]�#������Y���q�&�'t�VDT�*~qgmdԏ��Wt5�i�������y������z�����9�}
-�Q���e�ugW$轗~�C��'<��Cs=͞�w���\郵�������c���WPSj*ET�_�,���/����V��G
���M�x��V�����ʠM.�����>�V}����HM��,�L���ѹ�8���1���^������!�;���2����5b���i�~a-��yFG�G����#2\�P�,=�f0sj�
��}��* ���EM�F7E)��{}��4�H<��oX�>O~7Al���f��~N^N��a�
��+y�J�jaS��(��je�o��`
�4˟����.��D��:i�X�?O0���O�Ɨ"�%�S���(�	�"�*�U�_�#�̈́���U���u���9XV��Vm�7T�>sͺ%*���I�B{]j�rK������E<oa���As�!�o������1̥AС9x�^sE�tE��XC�f��rwL�#�y�6�{+!�"�ox	�&3~�)�"�ʞpLr��NI,G�;�[2O�	�7� �w`�23Hh�UZi��Fd����Y&�\Z�w�I����)�T9�{m����:�
��&<�@&�ԧ#�+΁�
xc�h��`Cs����|�E����Ab�>�=n�٩IB���#CQt����?<%�A��6�Mw�Ѳ�(�s	eH�^��W�}�@G?iA5~�ӥpO�L%�4����c/(���2a|ONk,��a����f�3B�W�`X�㮙,wܚ��WMR����]�t�_�4Y�6���T�Q�Oo�@�����,�^��䳷�r��ڼ:P�%�Ǽ��=��f^yLa���p0�#����i�����eG� ��Z"��C?�"l�C��c�uÝ�w[�<�%
�^\]4f�Ty��%�On�t�k^S��Yx���lS35x���1�+��j	l�7�W\�~�c.$f� d<L�|��±y��!g�c�d|~����}9�Ï�i�
�f����,�I���#���'�b������5�3ݶ�j�����0�x�w�9Eш�����e�g@�d�`������C]�Ң?���t�jB��7�Vw�N�����9Ew�"h���Q�iQQ��ɶS�;�ó	�Iu��J���mB�0(�'S�.|X��vȁR�rW˔�wN��5����~��Ǔe��\[��l���� �"%�_,S��tf�(��Yމ������|w?P�Q`���+�cJ��~��k�x|��搮�ƾ��u ^��H!�[:-.���2�T�l94}c�!�xi��8��f���w婮�]�"&��d�6��`7sJdU%��چ�̥�鳨E�K�<M�V���Δ�����;p��璙C'ǬΙu � �>�"�崯nNK����N�����}�hl��P��������ҶD]�a�tW�H�7�_��Z�,�K�拁��nR�b��E�Cm(�B�T~/ҭ3��D���*>�鞅%�օ��~�dh\�t��9O]Э����#O���C��(��I��C��?�'Xn�c����S\�}�����ϔwe���Yeu�dTXl���|fֺ����W�0�KH�#�\���?M#�k����i�����k1;i�n�O�]9��Z*^��G�ٶS6�{�H|(�ǍÆy3�ȡ"ͼ��bX5��J�`F���>��hI�R[��#��[�F���Y�7�2_���1�g9w.��0c��,�J8}�H�qS��D�j�ż�-u�J;	���0������c.�s���~	�D�!FZ�?խ'�l4��t���0;
�{$d!��B|���$n5�L��Cwn��9�d"��c���6�OU��Ԛ�GZ���jp֥��L��{�q�d&��2�uu�=��'P��M�C��F��/[�m�;��!���vt��LԱ:��}e�%��Ύl憡�Ys��p�l�q�BP�!d`�_|��B?��r>����A*�`Ǆڈ�ٶ��������F��.rM�pݝ�ǿ��&:6��Ϻ�Bޱ�_G���?_i�b��O;}[���nzs�a�߃A2��(�޽ݣB�4�IZ��v�vsQ߼�������:7T��-���P� ��ғ4I�]5P�Z����G&�-
�=�7}K\-�T�g�)"�������V��a�y�.��i�N�O���������d����x�4�Sg�^��Re�a�?p�)��V�c�Xs:��AP&� ��:�1aE���;�x봶������Sf�ݵ�_���r%yFkM2l���ni�l��$�F0�M�|�����c4��Gp/ �k�Sm�}\��]���3���Ob!
A��_�b�7�Yc�r�i���K��&V�> SU��o�r'h�\aŎ�$[��l�\.��XU�\�դ�	=6��-������q�\D&�����/NZ�z��VB4q�=�93�ZV���l�$�ȋ��/����a�<�`��e�>��d��W��a���b	�\9E��e�R�Bé	N��J�����,�O���zT�D%�����md� ﲅ��˗	k>+�;9����S��y�c�GA��W��$	�Ոk���DP�V��o��P:	O�&1@��MJ���H0r5�F���Mה�:=# wѭ2�˕d��lDi+�����i�b'�;���k��G>}����/��V,��"�Y}�ȫ��Σ���`�C�ǈ�`��*�ʸl��n` ����(��N�r�.M�t�Kq�v�xW𝂬���[�j.�?�zN\�8�\�8�O{I|;}�s���3�n]6>@��5����Cx���%&�_�"Wƚ8�2h���o8�2���<��[5���*�`�t:y���e6�<��ے�Ω&�5�5H�_ l����sG˛CUtHWMi�+���|�՚���0��S��N;F
�>�/	�}��Q�d Q�)�13͟��i��!�:�pH}��{���B�� <Wu�Fw	jk�(2�_���ӱ����T0ǧ$SQg2$`��_��ηK�;xv{��o���6"|��H���竪�G��<��mz~����dE��V��fl�cƕ3�\�1��Ûy\j:(6C�m�>)�L����0)���ʐ�	�����;�����"2��8��O�����I�\�9�j�={�����:)����xf���Wt��9\ ��,�D�\�F��p5nE��-ʺ}Ό�I^ �U�`�G�6�!�A�����$7��esu�j��aK���gQ��>:MU��Ew|řh��zV�I�Q��&�B���-Y20�D����tf|<���jr���:��w�pQ��F��G�𫅓��6hG�ǃ�B̌���MZ`�����^6��b�]��P��%<ϸ�	D��|K ә��)`�8���?/Qj�AO�������";2�*^�
�bw��HؽڇV����"zA�o �F�`)���d���fB�9f�޲t~��/{��oǽ41�[�����]v�����#��x���w�l�։o�a^R1,���2�u,�C�r��r�lz��Ts?)�S<*���s��q�zќp.;���)���f���I�aVS�QQBiO����!�ny�5s������M��&�@u4�g{�1�H ��b�ƥZ�b�e��y^��l+�'m�X�P_�����8���ô�م ]a�n����pzS`%g*H�+��w��b�Bu晓�\r����N���ܗ�5��Ĥf�{�[�e�u��G��_�ٌf<%a��x���eޒ�u�tV�ÉcJ���d�f%�qM���D�ͯ��J��փk��37��p�	t��Q�ĉ�(�`��,w���lB;�4���[�E������gT�?@n;�Q����¨��<��#:K{e��Q�hv)��]��ȳ���y7���uAMJX 4�6�	a��,�� ��cƋYύ�-�m��H��]|���?�,��5j�MT
\'N~�塺�\1�Σ��Σj�{-��M�O����P(�
�� د����q@H�Hˍ�h�=ş��],?��gR��Pc뿡��zy�E�<nR&>Nw�~j����;�]�7�.%3���IWǕPU������wnX��O-PI��CnUzj�/���J�~����ܟ�t��z�#|����5$M�#`#�C�-<w�ῴ��[��,qc�*���I�/(1 ����� �I�U�1X�7�'s�v�������&��|���\a��;�u�x
�R�����n����eay��Gf��`j�*���-�ڭ�u,p���z�I^�E�=���i���HzR;�#m������1�P���+O��wvo|�Ⱦޝp�'�j�K6�
d��դ�����!�f<뭈�n��z�8��bRE��6�c�\������_O{Ne>
�Mk.��?&g�i�9�i���
Ȑ�q��Ԉ�
�7ZW�ݛN�q�z-�60�+eC�S��eVC]��1���r�P{��i�X�g�"Gֿ�O��/��Bu1��h���W�/�f���.�?�r+�#|ז�����Q��Q�=�	�l�-�w%ϯ^X���&� �#����!��K�$
M�l03�{I��#)J�n<��ݷs������+[ 8f0�W���ޒ��0"�Y��=ۖ���f#��~C)��&�h���ˉ���$6�P)N@ m�z�V>���?���J@I�{���X���$�:qmY�tC�7Ңp_�Ұ�u³	f��|3��������}�皡 �[�\�"���K;�)N>�*T�C�`EU���I�a�@��7�!�q�М��En^�����o���ΞP;���a�WME����\���-J,T��[s �%���HT���Y��4G&O

+���6��1Qz�&m��+�Q~BS�7e6�/ R�<Q��l6>*ܲ�k_��)�[ʉ�c������
,~ձVYk�5�	7-8Bf�� v��u'N�U�u%���sy�2�Z��e�����vUY�]�H�lπՓ��V���[�"��^~�� "��P�rV=�B��(خ�]���>�8u�̼q\߃�u[-���q
�Y��μ�[�0�E܈'5������,R�W�}��4#Ҷ�LG��(�ũ�X��������(�����G� e$=��`ߵ�fk�SO�hy��W�樊G�7X����l���J�I��'̙�N�0���e�h����5#���&�m�I��
���0�)�>j���`�4K�����]چ�h�Dmd��s!�X^^�♏��۪8P�8�ǞA��J�
�H�B`��?:�O�J�+����g�٭vX:HM/�6LU�M�l�jV�{�QAz�oz�|�P��ն	,�K�`p��k��������'j���rX{����5]� �5�=�=���{�fП\[lO~�T�p����eQ&�u�,�-rh�(�.��ra��"�E�]UW鹔��_��x\ծ�<6c���X�ލAVҵ�""�P���p)l�������C�
ǝ�ǋ�
��fU���.5/�2�on���� D�����p}Xh��p������E�Wۙ��N��Ad��؝�6\����7�1�l���,�g��z��>B��
��h��ZN���{�k������y݌��I�M<��R]����I�%<}Z���0��՟K���x�uuޝ?igO�ϼ8��YH`,��tq�X�ַ~�]�>�aY�ځ����>G�[�\���P�AE�����.A0!�a;��ܣԮ�:�Gނ��ȉ���ri�Y�n��s��	�x-��M�pY��i�_f����+䚚E�1`��\�λ��d��V:�mA���[Ţ�l�Z� ��ʪ�Eܗ0�
b��u�D�JΦ��d���)�P�OO,����	�9�Hz<��f�|��Qf#B���t/��uz���D$~fh�^ɻ��%� KiR���©���@��>R�8?!���SA���ɬI�����Ņ����p����m���A_�>�҂�ǖt�&�#���A��z�x�	Ec�E��`#��H�R���&E��Guo���j;L��eG�ѩ�mǋl�g�R��q�8��
B���$Por_G� Q�Ë���[��{)l��[���Z������C3��YDd����D����>@����uքF<��n^�E��z�-�]�m#��dEP2�XaNQ	�i��F�{(�\v��]��bn��V����*�j;&��n�[p��`��&�Tz��|`$ve��x �I��Eـ�36X��r�'O�F�*%�U���Sdd�q�_�I��fT�_ӥ�M���Oc؞��w�]������?qpHC#���r���k����<�72��飋a�M�>�8��J �	6�m�죘d4y�$�����t�!�!F�S{q�`�2���R�iY��[̉~!�v�jX7U+��W����_rZ�7J�� A��AK5�:_������*p�l�Պ�v���>����u�;��r� �o�]ʧ&�0���0؆U �!�ʭn��:q�����Z����/)f+��7,���]O�iX�`�+c�fm\o��F�J�L���*�!n.5��T�ã�>U%'���PWMSI(�e�R��$R�qc�,`���;� VUr{?'+�dQ���/�Nl��H!�X�-�?,0�="=�xb�l�gpKҔ*i�"�ٜ'גVe��.�]'�-�R���޿0�.��έ�CP�����"}��i���90��g��ts��bj�����zh�*^7zU~��2I�P\�u,�cp��ta>���uL��D��BP��Ga%� ��a��LC�7J�<.���h��| ����(0�W:�<r;�s;ЍH�E������ݩ�Y{&K�����v���'��,�x�Ϫ	���@��"��=��K����JۍЅ/p�uN����I�N�g�| ����Jk� �t���0�=K2��pр�<��W�8�*'�~�7H�Qi
Y�6���@��5xa,d��?�[ʣj^�OE�].���f���_�T ��X}b����x��y$+����2
�b$%��Ŋ{�a;�P�'��`���c����h��P )i��Be�$�|�J �]0M�P�d
2�E b�	c.�_���սiP̑�G:4c�K��u�����.�q{�XrM�H���R�=�5g�{3��&��Bh_3�,�u���-�Rݚ�����DA�;Q׬oZ�%W!�s��
zƣ�X�r�2�H��ط�L�O$-;��+��wݱ9��Aš�3��H�Ľ�*���j�U4{���N�>��Bj�[[@{��P��H;	I$%%!��~ʃ����9�Rn
��Yiv��Y�7�N��{�F5���������b׶� �W8�����3�y�
3F^����l^�и�2�%O	�$�
+9{`-�U=,�Z��d�>)�Q���Oq�;-�����-w<����4Q�_˜�,H�j �sapZ��@ ��M����	V=`{Ui �q�.������>����:��^�~ܚM������_S�|��$2�q��l�C���q?U��ߢ����/=���\�VJ�U����|��6�[������D�hL�Z�tE4Zc������o�N7�.���X堫M�.�7󰾍	j����h�R�}�]�U+g}%p�=�u�a�n4��9��\�`}-5�ґ�����4]�a"]���a{����\A�G5�����m���Y�C�?�m��G
́!��������H$���W̎&6�� ݲ���l�+e7Qsc53�yR"ɒ��ѩ:��([�,H��e������+ً�c�oȂ�;����j��_�+P��i�B0�X�|��[����F6M��#dځ�P)�2:�9KV��S��޻і ]�0����m9��Z�2�v�%����2�L=>�?��,�W��׸�d�-�0v� ��R�ȶ]�͜ ��&�B�4L�X~Ͱ�Ԕ��h��o���r�ZD3]"�X��|��s�5����fjVy5�08j#�Q��ǆX1����3b<k=��.�=��G���ulM��ӴZ??y���h^p����~
Hߘ�+���:�aU&����e�wn��@�Q�9<S��y�P�e�Ǩ�p	u��r���#��w��8�U��[���L|������	�ڠm��|�p(��c�Z�����4rf���{��r.g�*B��m�|4��8#c�z��>��+��2n��߷��]�`X��o�R_`�*B#͏_P��hG����U���j�q�8r��k��Iz��<�E�P�f���qW�� �3 5o���[�7��������K��jrBhZ�-�H	���y��[�|:���� B�cP�1{+e���*��G�;�>9�1f��;�'���&Z�g�ݒ?Up�^� K��`���i m����Aظ%"�)=��5�Lti[���R�'�x�"�л��'OR�粖��@�t��</L>��Ih��%��<���ź׶07!SG�����R��p�H¬_H	}�/��"D�����d��
�B�]�T(��j?�I~�&�1*<J�F5}ʙ�k����k��LIGOAn�i0��W�R����2Lp�o�(���z%��aL4A,P� ���&���϶$��\�K� I��pJN8�(��X�p�b�W|�%:�mZ�ep�&p��ZC����q�Ӻ���p��:ٱb������Hl����w�?>����L����|˦�?�6X�T�q���	���p:͜���:Ŋ��j�_�\�,S�~D3�m��Ɇ�U;`�k>.����i�>���ؤ�'��0���CTY�:�D�e�#Y�h$ �j��GY8(���<�@�ǫU%�H��e���0)�����kh>:e)��}:���I����"��j����"�ތLmK���`���C�B
��,�x~��7��:��#aw�<�����%,��\w[�wv_��ɣi��i�Ԡ�i>9MFP�W 
����Ձ9X(�1N�u�3K��n�xh@�  O]q�-��P�FVw���s���"p����[7l��b��3F������o�� 	tc������ԇ��hb�Õ������+q%wDL�dF�꟬��N�:�Ң��Eu_J�#I\������Ր�}Vg��g�u ]Py\��؟�,v�?�pA�]��q�4�x�H��"��²`��c�́�DtH�H�������?�� ��ްGo*����j	O!�3���c���>�tYiN�LٙV�L�r�h�ll����H�A�v;*�ei��f���͞�G��	�"��}n��F�I��x��`u�"e^����#�S,\��i����d#�L�&G�M�} ���_Y�~=���S���xS��v��x$�d���F� k�H��|#����������G�`�����O2z�߿g�\^��ĸ����[u_j�6������:��[�4�ݸ_��ev[hD�P�#="S;t�|�K�)!��l�D�'�'��c���|���!*��UQ����A
;l��[��\շ�:荄�ۄTH��]!� ����)��"j��\L�V�m�@=N[/��v���Dn����M�uxN�{n��9c��&��L�mP�c���B�$-6g�N�� �k��b�-M������k�ZY���:��Q�Ơ/�-/I��H6�*{�M�H�۝񷉦���>��$���F��* �躇���<��[��ϝ)I�S��,}C������l	�@����:{�:�J����L����$8��%q���4��Z��G]�w��ݽ��a�a&��b��B^�H(�7�$�LnA�%t�\���?�a�������X�qD�<oX���L���F�3uȊ9H����V
��������0��u�~S�:��|0�8#n�so��;��og �tC%Yuy�Ģ#� _;Q*����~e��3J<�i|HT�.�Ci����L���ߗ$s���9T�[�[�+�)턐��^�e8��{G �j�(o�u�_�ش��/�(DL�Y���W_O(m򬡅(=t[�+ ̃�L�M��J�YBx��!�-4R���^x7�"�)�=h�ŵ�Q_�us��Z��L�p,2l�g�9��B��C�"��>�Մ�<��;�@"�_���9TO�>|�t���l�y���ݡϷ�O��B�ck����(�r#Zv[���L��mq��}�����q����=�()��l�__����P�%��so��ߴoo�%�1Qi���'��c��dF�c�����ήr�{�O:5�e�4ib$~�EkO~T�h��<`�FݖV��U������ߴ��ix2g��n���;���!�F,^��o_�l�Y�@�|Ds�_7���ӧ(��'���ѿ��G�Q&���~_���4J�C�ڕ��e<Y�<E�_��|�/+'u���J6z0*�U����	6ǿ��]Y]����#�Tϛ��"�G�Y�w��'B���8����Թ��V��]�J7�^qz�������)�c�Ԉ$�Ow8����o�1{��$�d�l��K��_��K�^�~�6Mb4�[��F��̏�R�s�	��ɺ�Ӡ�\���3�[�ȃ�>�I���qGT �~I�.��p��K���$C�r9�=O�!��K��r`}��wR����,�����#����H&�L�4��a��.6M�sFG��ք�9�Ff���x	��_U�N0��B�$V#��<����Kl9Rj�����Xyq�A���R(�zV�
x��Z+�^"Qgm��!Ax�e�}V�m����~�
�tk0"�K�o��Ϟ�ޣ�٢�-�L�
x<����;�Wib��ʀ�W"��y���h��HW#�@���jP�!��76'����1EW��S�m�n��Qk��[C�]T��Y��֫�x��w���1\G<Ȗ�%�^���R�&���.E���l���/�}+�گ�?Ce(��o� ��� j@�U-(3�`��P`������R�)+�Y�} �`�����X��o��q�m��l%��}��q\��E>��)�@�{!l�?��U`�]��n���+��z�oY	<kƀz֞����V*���>����\?QegjY��!^Ñx9��5�c{����;x�'�S��82kO<�dM	��Z-�PUå1�U�����5�k��(hʤ��]�W�y�<3� 5�	�5��.�c <�1<��5�9Tmx1-���(���]ic��. ����N�Iǌ�p"��4W�BR�O��^�g�epʰ��~�	��e�����uY�
�x=�"�ta�iV-���1毻c�:��jT��sv�ƙH$G�e�{ȳ�?�����.�?�エ�>D����0^~�J�d/�1��d�c�	_�̴�~���ν��n��[[�,�A�O��g�}���O�9U���&�������)Y/����\&�Ե�^�S��j�Px i�!i<�
J�6�}��d�*M�2B�43+o�L���fߗ���m�U1�ێ��
N'�'�M��ի����W�jV���t�������d�|����/���8��I��x�*��P6+������E�wXK��#��,������@��_�Ϻ�=$=�~�� #�t�-�#}�Og��&:lQ��k<h��KMw6�促1�-�{��WO\ �h��dy`#\�ՙC��(�`Ҩx���۽��#i^�*\��Դ+Oc!��1�.����E��&��\�R�{�N�-Y��\{PJ�2��ʬ	�tb4��L�)MŹ�OS�ing��l�����J�js�Bh�]dڕ���b+A`"|Pf�*���kzg�Gi*��ٵ��d`އ �o䎡�Q�Ղ�bׇ�9$�/DG��~�4N3���)|\P!B�6ҁc,�в[��MǨQ`�ǝ���ٙ�jE�9�\y��k=���K��Xp��o��5�s�TXL0�WT�OZ��.&��j�����(��{�h^½��x��1��-�]�KX�́�U ?Ӛ1���Zʰ;� ����a�[܅D7(Qc#�X�c(����;y.��ç��V��%���4���ae�{����@<�H�}v|�L%d�f��\�� ��R{�jh�t���j�k��݈����}P��#��s�1��U�5��>V�j@|k����h��ʰ�v#i�GR��Z��ԝ�7����g"W�`����O?�8��j���S�J�i���%����p����=>&� �@�C֓�4JW�ĢBW�����>�)���[��`��>\5�ݛ42\�[M�SRVOp��v�?�r��ʌ����"V��� ���3֗J���#DF�v�����ؘ�+�nS6V0N����M��.�_?_��p�G4Ń/.��a�e|�D��2�>|�-�e�*ހ}�qc�p{p\;�����=y�Bz�W��޸��vٹ��Hv�I3����N7�U6
�RM��Њ��AzQ��˰]]��x<�i.����ÙƗtPo�H���_<�
��â��t�����qi,�)�$O�c�� [W��T|�	���2 j����wd%��C�ķ�P�����Y���A�x9�OY�Q,`Y��4f+9C ���C)���<G�������|k��B&���'w�J�@���w��Bߪ��*~ Z!|��+9ťc�[E���`�'�'K3�Y{��v���.O�{��;S��j怞���d��&
���xM�>�|F�#�IC6��b��ФQ ��'eUS|Q�KIu���o�6�+i��	Eآ��n���W`T�ug�z�����ƀ���$�Y�)O8�_EoKX����0��S�a�^���qM,����H�x��g�^b5���/*=�3�ݡ?L��G���?�S�0�;/4|}�8�b	�bO���aW�!< �N����E��`��َ[	x�,$^ 4�m���K�x�!; ���ni֮� �%#����ܹ"�q[r���Zr��%kY�*�Ԝ��,��
_��i�G'�F�a�����g�G8����C�kV,�	X����,�O�LE���]�$�<D4^�<�u���<aYS�E5n�7���=�'�zo�,����F�>W4 &����R�N�N�R/�@�wa
c��b]R*!2!��ԟ��{&�Iv����'k�Ƴ���YH���+!�+2�"Ȝ0M��k��8�/8��#��i�����j"TF�H%i�~��Kk��5�˽[gPk�X����.J�Y;ymQ�
8[U�o��Km����C�f�e��g�mc�^⪼���C�r�����,ٌ
��&�x>���	��F;{�qK�g',�<��5���D%]��>����GEH�,�S����+�9�/�Z�c�����LNb?f�u��뫜R	+����a���BZ�>�u���큡�e��?��eSK��|������@�(~���	�*&+1����G��y���O���zr�P2yĒ�!�S��i1 SL�=;R�L��=�*� M�d�x��^޺1�%C�	�7����'���˃��2���ډ�O�� �k�W�����-���Ӷq��x�ky����N�{�e +�BK�Tˬ� ��X��뺊�ϑZ���Pe=�W�\��p
^���F]aL1�׉�1���6ζ�RsS�JZ�Tu�h���c�MZ��p`�}5�9�:{�@N}οK�,��~���T�T�=�ٹ����2 �FC����u�����n�J̮Roz���<@K��"��� �㯱ۢ݉���Ob�>ŋ��!��FG�+A��/�u���w7׏��r�{��D3�c�ޜ5��t�'�;{T���#2�i��-�{�خ���2�2����u��-���(?�(�<��n}ǻqؑ,w;��2q��l��&���vժ�G��Fī�$^�v����YA��	��d%_&cCg�����g����]k���v�OW[d3P�0�.��֜"����6�/�\�s����魾,-�f��I
]�y����a����$堅����I?eH"g(u�-c��b��"^6̠��M�M���ca��X�<���k�;����-�{�&�����<���H�szn�(e;9v!���o�y�'��h�C9m��/��T��{}�"9p��z��Ǎ'�s��@��5�W�4٦7�W�^@�zs��^�* hx:�).�����_�!)��q�����<I��f.�.j����D��A�5z���K�>��}�,.eB0J���g�0�~��J�PQlL��[��8����|�����Ǘ]a"}�ё��S�
f��4�U������X�h�E�(��5,"�%C��ec�
f�K}�j�V�z��"HO7�M�]c�ru��z�n7J�n>�lbD�����]i�5�Ǩ�&�j��"�?A�R7_�@�P���,�D��o�����%G|������O�/(�m��Ӥ7!�e^��/��gsE�����.�v��� S��,���b�9�FxMqn,is �K��3������E+0�˝�B��U�"?B��&�L�V|Wf�ɾ_Q@���H�>L;�F+����"����5l��^�ʤ�[��2� �j���i��K7I�8;�G%�����E0m�����v��;evdn}x5A�~�eސ*j���Dm�DMf�
����8U#��W�צ�dhXR�
=Aǆ{���\>��Z�І7�lZ�����&h���Z�,M��S0h6�V�e�>I9J��Au����-�@I��A�Drm�A?���2%|���`�N�d��=���V DC�`-pD܁��:��Z��@��*kwm����|��m�:�{��7$�X�ģr"�S�Ͷ2uF�43����?�N���'F��{�8��vT�Ͱ�Icg��@B�L[*��ǘ���$��uZ"y���~�b!Цc������g�'��8��[�B��N>'�J�"*����Ƴ��x׌���
����<n��V�������R�	���L���sY8�M;k�c{95�8��W�V��H� Q��2��Wײ�b\4!����ݹ5/�m֌�CK�1~?�����|�����u�_�]tF��'Hy[j��~sO6p��-+H�F+��������fW�� XU�O��$�#��VAI�TH%4a>�u|�`Tf@�/as*����Q��hm�[)
sz"�g�w�בn-8��4�s�o�X�M�pR�~��w!�_ �	��zj��y���L.y�}���Q��C6��2Z$�eЌ��V_���o?W>�����t��R�Z��!,�������c��B~5���h�[��l���qL ����­4N}r��Շ�(Y	����8h.F%K
���ɢ=���+g��j�P�3�Y*w�_4�pȬSEL�%�y�$R|���Tl��?�����#�`j̇O���?�; 3:EO{�NQh���\+T��N��r�ץu���7,��3G	؈���<��`2��*/&�����aW
�d�5��,wc��̾CY������P?/5i�U�m$���X�p�d�(�P��~����T��� d�
<�瘵�oc�[�"/��^�qJ��[Nh>�n�iYW7��)Zs���X�	�Skuk$�Jm!4�b�F���Bbj�'�:lΊBv����N
t�����=@��^j���Š��۴���]6ߋB6fl,�����o�e�IC|׋��Ԩ�Q@,"
�';��T�	��d'<]0�L��Y�9�xje�'�����Ovώ���M^J{�*[SӼ�X[;���Ҧ6>2�n�쬞��� �?��� �I�3�8S�H,]�%�j��������q��K)l����m�C%�q͗�vڝ��b*�_8�����FwU�_���+e���SB�}�y����Z�$��x���îG �6�3�d�GNBěeNݚ�����J�Wa7-|˜�� B ��{�f� W|?���j`��0"�`��%c��6ےުc�+�?'l������REu*Y1���AI7�H��qi��6:P�>}��Oj�	��<��ԥ���V�,�B4?�2���J��U���[L��"���X-b{'H��(����M�3$(eI=�g��I�O�dB��k��E�E���,R���Pj�D@��${a���b> n-�{P�˽���ј��B�|�S�-�Qb�'�@��@��f>/��H�P��S��HU��[��I1յ�<��$��E�yi^� �͸��t�#чg�I	��\�y�����#�:�"c0g�c��������B��hӰ�=����n.����vڕ)������ ��i�I޽�щ}�%M���9�@��X,:ps@:jC[0�#��&$�e^���7�
X�g��>ꩣ�����T��W����.��U����e7{4�+�	���)E��2o�^���znb��ƌ�wt�Nx<mڠH�S憌o	����� �U�����'��0�x�k%Y%��.8݁�q��"��웓5����E����eq����Xj=]���j5�D`���li��3�W���ٕ���m�Y}1��Ú�0�p�ێ��O�`���:�z�����T{��*��b�ߊ�9HL��$1����_�YeS�Kb����Q�A�]���іG �`.YZydɉX�Px�m���+�}�Θ��R���$Z����'[N�����f�Xh�������Iyc/ �i�b��52�DuO� ������E���C��h�l�;B`�*�ʷ����Oe�ڻp�9�n։��v����GTSVPnc7d����������]XE����)��%�6��@�Xq�QVs�+5��ݳ ��
'�ՄZ���U���F9���k��1�� v9q��?��^���u�i ���NTM&�pB��t���f��r=�}�-=e��M�	�0B��qA G2L2%��|u��C����uI[�;y�u�з�>f��(i���3կ�m(G�q&i ~���-�_���CWp
S{[y��0Wq�6m�#��8u�X��e���I/���֣�#Y�T������(H�J�1M�G-|h�����a�<5���mX�|Ձ�$��q (Z��W�F�b���9�'�y�r �rM�Qv�7��x�0F�*��|ҍ�&L<L��S8��E��&׉����h�RT�����O�b�ȧ�D�X.��U�t���a�	wπu��N�aj�i��؏�QફǼ� \iNі�fQͺ�s/R����,ܺ�� |�C��4EE�����#:P�4x�ۨ~�LK �J�$M��8��O@����tc�X��#�%���];�Z1��Q0��c�*d&��$�oˎ��J
�m��%��0ڂ��	
�JY����K3��݉�sS�����%@~��O͋���ʔ���!�����q��OG���q��#�d�gE�R� �����zv}��[���'�>}���2��GK�>�3�5Ww&m���,�IةT�C�`zZrݖ�R�R��L�f]k���P���hG9�~�0 �衳�1�&]�X�Ҳ$��C���h(k���H�[=��k[T=�;l���n_�	� ��u��I��;��m�������d��99�-Z�W��N9��h����}q'$����F�N`�O�1g�W���W�b��HL(H}���H��Z�3��p�1b	�:�(����/=<��s�y|�tB�(C��o��f�>�0��mX:�فKI�R��-_��:��T�2�qy.���h����3\��F��:ʂ�sD�����Bj�g��GO�����:ci���F�*F�]D�D4n�8e�NF�F�����2H��Z�z�c�m�g��/$�Xй!�0��FkqF
�{�)���`pw����+�ԗI�1�,���#�칖[o��iߴ��C�j���;F=�����-q��
'+G&Ǔ8 lޣ똢	�������.�(qp�Hϓ!��Y��
��h��ɕlegBcem�Y^���&Ũ���0��Kw�#6/�p����zN�*]o��#�>�q��������Pm�7����A�&�G6F�K�X\K��IsL��(�Ȃ�b��~���^6�r�F<#؎����9����fН���.=
��髻�쐔����V_�9dA�f�h�p�tc�MZ�!�r����fE��qpw��5����x��cY���1f�3��:���p����)�p�m���j>���Pg���Poa�Y�� s	�2��k�K�%�n$~��F���Z8&��Ⱥ����Գ
 U�UkHe�6��������$��$��_  �g[�8���`9*�G�`i���<�\�BԴX����>�nk���Yd� ��6�pwZ#�C�#�X���A:o�C@C�����:z�S�М��!�Rq��\�/�� �0�����g,�����.ՄDA��m�h��c㨗o���g���6��e��0��F��ς��u�	K��qH\�3-��LN/��i�dmF�S��4uMw��)_a��W�;'�`4����7��'@/ew�������@��Em�������7O�F[�5�.�X.?�:�t�~��9�����Ox��^/�a7ا=�&5��B�9��6��� &"ٲ�_�~)Լ%L�WT�$YA,݆�|1�VR��-�\Eq)|w��I��,T�':+s�������.��p���=o�jU��)��t�@���A]Z4*O��X���Ԡ%�omj�d��4m���̐i�[���i1a	:��Z��i�7��ڹ�o�؇(�+6�7�O_��:��ݯռ�EB�R+rd�?�Ċ�.U�j�C6�L��b�}���d	&`�������բ�1�ܳ.�{��&L:�f��n�=�`�ѱ~K�dAa��i�Ƭ}��pQJŗ�x�dAM$`�����t�K�r���m~jQf�0��B>�
��y����v�LvT��쬾����mbi�w����Öf�X�{��ħ��5-�	�7���Ÿd�N�%�j�Xi��{��w�.8�뒿�-3o�aY;qm�'ܫ������ �*͖�+�+q�bb�ޚ$UL�'W�H �jr�丐A�z8��Mj�����m&A� KC=���]��� >�7߉A� n��X<� �'l�5�g]H���?�A|&�q='r~�KQd-p�s����Ph����>D,����55���M_�r�{���'{zj��P1@uƱ�_�|�E�f�d�c.���{_�N��	؎ޖ���ۈzn�����ͩo��':������}�L7�8�S&I&Xi��8�\���kO??�~��T���Vt����N7P�hm��s�a�vJ��{$d\}=�V�������fZ��G�m6��K�i��W�}$�%� ^,��S^�vA�x=и3>�"��!���Σ��}�*��������J��_r	�C_���(��#1�Ͳ�o�����.IY��p��0���kR�i�Bf� ����o��FA3�K������ם���@9�XS�*�M5��2��4����n�^&*������`j~�Rm����h	���	�9�oT@2I�?[��Q厕D��O%��"�"��#�D�WAX����o�o k!� \�M!���{K��� � ��<X�5�R�B�B*��Լ���cÖY�v�XT�#y�S=Ql��80�? �;�#?x������u����R�VsG�����1�B�K>쫬n7U�|�*����}��O���,B�+..�p��G�,m���LT	�i
��w���9���h��Q~���x�����0w�:ᒬ��OȮ��������Y�Ȉ�i�$Z��nz+ͻ��>��Hr��C�^�W�F5P��P�D̹�·���h:����a{�|�Bi.�����^s�qiS�s$:���*[�L-�e���-�W%*'�ޯ��-��9�/j���d�ނI��8�2i,Ú��ŝ��YF�b���y���%����Ԃ�HQ�`V�!���!I^�K��PW�$�2�%�C\� �Wz�s�xz����{\
��YW	
���5w[ R�~!�[wn���Cky����UO\�v��;'K����=��(/fCN�߅u���gp܉��3CG�7�4;_9�|mP<=��F�e?���	�`����qʗ<��$�k�����!�ݔ-h������%c=�)�3��r�\�BKw?X.�I8����|s�V�Iǉߟf���Acל}��"��S��C�˂�c�<���KW�W:Q����f�I�C��T����w���0rcƞ?\�uG����]A��7������Ҽ���	Z4,*�x�$3�����j`���3���ka���.�J��_c��
{A�5�d�����s�y~��z���❓� ��oS:��u�+e�j����D�x_L`־y�'L��%~��늴E�S����Xe}��t�1q4�(���c�B�ߛ���E�7���1=���L�[�4��|�]E����7�D��ujj�cu�tI-�ڌ����Z���G��VJ�(9�����`,t96�>�Ƕ-Z�=���D��	ƭ�fs8rr�􀃸�Ӭ��Ơ���g#:����Xv=�f���nwx�*�]Mq����t���a1ɒ	b���:��s�8�ރ���+��cs���,��c�����?Iu�|���$`��c/���q�&�~5R�_�J��"��Ǉ�7�XLV�Q��")3�'�*^ׅ��lx^Y�o֝	TP�ZjH'�^�3 �6�R�R1+��4�lI� ��U�K�Jw��tb6��8{i!�L��j������3�T���"Yǝ��^�[��䑦�sN���E��J�g%���7�dE�e�9�)��?F�B_�n�#��&$�l5CX�j.\��F���I�2�<4�?�	� ���]�Ț���R�n���.�b�Tc-��h�w�IQ���,,ד՘�%��ޱO!W�g������ek��*oE#�4�_� �#]�N�դD�50�.�7.�ġ�On�Ǜ�� ̼�S��&�6-��l�no���^� �}	T
U�> �_.U*~Qz��´��b�b��~l?�F�7�B�o�8A�0�`gJ/�5˭4�d�@x���0��� �k��3[�0�׻������M����5�����d7>۔3R�1��VJ�U��u����!&�./̋
�������_9�Vh9觥	�nҩ�+�0H;���MI�Tt*��@7�3d��0\]u�uQ�1~��R8�p��w�:�^�ϙ�94s������־{�L������*	TdTt�LY�x�Κ�î��Ë���M!*N�P-M�/��{��/yEKY7�8e�ٟ�hX�������7φ+�4gG��L>�jԳ�/���G�eM%J>��p� ��0���U50x�%���i"�w�K�Q�7��&_R7
�?-a���h6��_<����������2��8ןG^Q��	/Ǣjhd9����V�ZF�F?���0�a�j�܋g�M��q ���ᔩ��6�-�a��O#Dqܦ +�,������ m�=��`��"�Vw�SzDf�_�\kr���r\�a���]��"��2<��Sr�?v���W�󽑻c��P���S��r��l��I�旋Hd��6K�U��=!L��#\F�0�(Sr�bFmzDF%��W0�4�WMh��\�N=���2����Ύ_;�+;�������(���8T0oт��MB��6L4�F���IGe�U@&�8�.�ļ��Æ��$5v;��$�ˠ�Bձ5��Q�hE�b���D��u' �%OPX)�Ą� ��v�i�z/�F6.�}����
w4�`�Z�0�p1 l0�*h���l�����P?W�X���RI�QsD$�p=�-J��@G(���M\�� ��,� ��JC�})6�G���/�^Vmr�iF���CW�37�E$�}"	���`C)jt�'ޘ�L��B��}��p�U]�ء�J�׉�FJ-��P�J��z<�K��k�%v���p7�̜��k��국\��qGe�ݲ�T��� ]��Ն��N\D��o�k�vT�Κ҈k��ԑ�
0�W����W�s��� ��?�I+�[2�/�i�R2�=^8��sXo.��E�9��9�j^�M�M���ы�Ra� ����
����U'�$Fy�AV�O��%���kLUw�V�<ܾ�^��j:��"�hѐ��3�.^�}�z��p��_����v���ulkY��1�5dӟV6�`[�=1~|Ñ�X.��N���)�;��|���9𝞷��Q��wq��~bn��_BQ5tſ�J��q��W��9�����L%
��i������聣���M �W� �G!N��~\���P���*��O�����s��?���<������N"�[X���<f��w7�ߕr� ȧ�"�p&}�����j� �tr����G�Y
O�t�����l�,3^�H~I�Qz��$z�-
G׷ӿ��D���[�|5�-�Ѱ]%�:�9ե�b����?:@WC�ߦ~p�ضi���7&��`����,?͹���cMȠ�֕���O��F�QU�؏�::�P��y؆�y��xȭs�,�&�	�A�#���7�]>O�{#��C �ps�c���5Q��
��_�5��ɫ��ph�����I�-a�vץcC����߹��{�ય��f���ˑ���	���ӈK�@|��0S"n��<t��O����������(_�])�[Y�J�r��}���w5=Z�T*����5��)sО{t�Ο�=Y��GY s����֐�9\��Plh�aT�S��\k��h-sf^�c��e�6)Қ䵺N��T�e���NA�C���z����yB~!cܫ��}�ҟ�~�E�h����zl�CB����Ծ��ɞ�c��yU�!�b�
 A��H�����1�@>��P�M3国�^M��Od�Y�)��b�p�x�$i>aO2%��;�������pj���7R�*�*e���J/��b���=6��@�o�QD#f�r�RL'�cK�T� �9�8������Y=�Z����խ�9�a�a_�#3V,1(�
2Dn���/���&��r`$�!+�
�?�R�4\�ڨ��(�;��"���_f��]]+o�҅� 8�\­͋�fs�k+38΃T7񭣻�P6~C` S�^1D2i����R��\�����|���i�X:T��d�&}m���ۍr��+eP$�g)�B���Ԝ8��� �&�:�d[d`?@#�Ҩd� x���l8L������*1b:�S*i�Ю�}mI��#��	�CafB;h7��'���P�o��B�����S4I�X��=:4�S�����c��`+#��k���C+g���< ��ލ9V�X�9��ذ#�2�O��b�.�R��4]V�2ݮ*������g��P��BK����g������n���܇��ɘQ��ʅӀɦ�N�N�D�!�*�1��d��̝ذ�-���p�	�
�R��鉅�&Íb��������Џ�U��F�r#�=s�E%W��z�[�n����=�'
Sήތ��_�r�2#\pw.)�A�.�NX�έ��"9��#��gk��Or������ܹ�j�A�N��R#H���y ��ܵ_�ҁ=e���BB6����D���($���P0 ���b�Qէ���Cn�;�,��j2��F���N�� :�s|��W�*�	n�;K���p�q�08��.	�8�2�r��O��$IO�,�Ih=��ѢAj�Mݤ�z������-�t7$e0&쿱�R�?��֘����Z|��%�W���g�m4E�M�\��Ե"ʢզ>��m�?Yx8��Q��5��:5v��"uTHx�1"�ʶ0u&܏�J�eGJ^���&W�p�����Q�dP���esvS7o��w(Y�,$sA}���Y#�_�#��5 =[s�`���1M��t���������/zw��m]:g�Ni�R ���`'XN�ni).���9�� ���I"�eF���������f���!I�&����s8JVߒt���Aڀ�A�VP��-���pLa�6?���x�F+��OF5�<�8���:��W3?��QM�pktsl�g�qTB�������9��ϴp�t���8���i�hܟL��k�;d&Y/�9��>�)�ho|/�c�|%PG�d���\ j  \�ĺ���Z%s{ha�C��ٕ�g�-���;�2��)fv�֢Iܶ&C�?�)�>��Y$Y5a���a�8�4z*�߆�c�!]Iea*;p���vӔ�����8�x �&[e�~��޻���qpZ�`ԧ���sO�����y�m(:+VhXx�S�f꽕]%o���ejb����_��X��JS���ϘVO N��^||pg�=�4���\�j0Iѿv��伤�qN<|EI�@X�������#�2Ͳ}8oX�sY�R@�^��#�H ��`�嫤����ʢ9�K\��+��Qd�F8�����b��q���"�YŞK���K�%�V��򹥔FD�=��Q��p43��B��"��q��+�ݕ-����p�]3]Ma
PV4�f���}yDlh}s��W!���mi�Nh�1װ�J7��V�z${3y�W�DUg�W��6V<�;����r�>��H*�;����$�[���_F�e
;�mEq�$����Y�'������l�h�i�"�j�C�^$K�m_��2yn|Q��$p�&!ɐ2�;7z����tqjC,h����\hˈ�eݪ�BC����r U_��'�=�R�AD)�N���C1{�fF<�e�� "9�\��*y���j�y��m����*�@��o�B[a��7���q'�,�L����U�O`��q^�-{��Ǜ*�Z��0`�j~�F^4yɸ��՗��:ư$ѫud�wJ0N��r�L"��7NX���O�a̝�S� q.��=���S��%Y�N����&y|a�s����-?qFݟz�N�1��;�jh��F�튉�
L����xF=�w���/�4�f7��I�Eu�t%�M�g�_���ߐw�!�p�|t˿��LũI�H���>�W�i��c1�\�A��b�àp��HՑo���&��߱�U;F����r;��ۮ&NTFđ��cs��{dMI�/ �0g��e�B�F�g�؄g�Gsq�=`&>[��!.�^�n �a���q�pA���-�["d���1f��S嵟�>"�%�֪��Z�W13a�.�޹�g7�/1f0i+�A�T!ۏ�q	�z_�}3e���U0�o_��x)$�Pl�{��mh�k�Q���4�l�D7ܥ���<��
s�Jc�sgJ0�(Ps�*��c��k�v��Q� 0G�|>ڷ� S<�.��T�8ʳ��Z��'�J!�D�.�￱TQ/��������*Hu�7�r���ӄ�fp���>�|^�R\��5Y���o�0�J��d��K)EW2jD������s�� =�&>ۯ�ۺUo���-��(�po2�t9r�~
�C%�����*�1��"�"y-���jKAd&8��o��g��h��ˮ�@+�Ц��#�'y
F�)8GJ=.}���>f���;��I!���&�C�ǥ�W	�� ��5�-��zD�-'�bT9G[�� A��%,��e����~Q��)�#g4�%�3�=УAn��M׉�C`�m�>��驩#�g�IJ�V[�"Z�D!f�X�
�u�����y�u+Q���KǑ���7������st�"
m�F�vC�q������x|9I}?)�s�-�"���(���	[�(��w93_#�iWJu'Rĉ��h���	����źj:?V�������5�(�~�c��I�!��<���R�,|�kK��Tl��gb��Q��̋/r �9����k׿%��2b/`�����I��(C?m��=�w֙�W�8%����STTӐ=l,�ȅ:�^b�f^��	����F�O�,��%n��h���U�WH�C'{��tQ�L��p-��������M�)��w"@�-3�MR3d �]
A_'3�����B�d݆Aa�H*h��AIJ��3�71�J�s�r��%���U<�Rm�Máٯ���Љ�{^ew�dD~���W �9���V�K�=�1��-�5�E��쀏=�������َ��K�#�H6K�X.>*��-���C�&�lA����]m�!�mBԚk��rA��uS�/�G��Lq@��2EC4�1
����5��i�K����| ��
�o9��Z���-���Y���$W2�� $kpv�3 �ŖĲ8<������ Ȗ�$@{]���+&�Rj����5�8A^m�����֔*������#�m�Z�X��($�&�*-���[ 8^o��a�� ��R5�kb�['�����c� X8�T����O1���l�8��L�p��u�^.0e��Dʪ:�#��P�"c.Y���Si��dm��]�i����.�R��d}��4����7�\���J��z����	6n!d]���
)Pz����/�����Z�'�%$��ęIr�+]�dΣn�H���R��:��?M�]�:����_�X6V�x������' ��i��RD+��Y���A��`)�mA�׭&,H�pq��Բ�'�":�e�������1cXY���K���X��	}�b�&��,���j\6�Y���/kf���ZL]�6Ky��fUU1�ϵ�U�������,s��4N��x�z�.`���ɻ��/�2�����GcAL�ܽ*'�3�q�Kq�#07��ZVv�����@�l�7q��,��<y�I&K�;�u�7$9�����A�u@Qט�ܲ����p���j�Ɵ�z�YYmq��ȸ�����`LX>"z�+h�W�!�{*8�A��M]��Ey�%��w��rTA�9=>*o;�y���=�����6`���U�6c4`F���T�������Xo�������6j�� c�����
˲Z�]Z��G�H�$����Q U�v�2X+!��:�-�$��ΦX��拀��HE���鷙^PG��(�9q��T[�[B�@���e%����uL���wk�mg�,۸B�wvX_	v����J��oѨĞ��T�󙵋�6&��_�էYf)�u�#]G���0���N
�z4�`�{��L�5+��1�P:���ȡ�����5�L�O�	�j�
�Q'p܂[RJ��k�ԉYC���L#�����G���gÓc^A_n�Q߅V��������{4M�����F�� wi
'5�E��h�z�
��Xt��xs�Sv!ؼ�/��J��~�VZ��m\�N�T��4���:�YK-27��7��}ׁ�"%�/�_nGम�HV�鍪k���r��K.�� dU,Y�R�E���`����d:�t�g����FO��	(��܎.iq�7}�r�fz�HB�]��|F�;>�D��? �U<1#o	��E��Ҷ. �HL���9��|q���z�J��Xci8�|iS�h��_��F�_�o�v�l�����	g��H�fI��]m�"4��	5�Ga��a�8VY`�A٘(�y�z�*����=G7��Q����%J�o�.�kD��?���R*�ŝ�X0��%"JM�o��s��t��
�dэt��-L�U1�����z[K^��ƌG_�C1z���_�~s�#��.��OԨ�U����W?�	�/t�|�.BA��fĈQ��有�]d���{w���:��Yvwn�����ϘSO�W3��6��^[�����댼A�	dk{(�M�@��v�忷@�+�37C�ﶆ��c#�d���[z��sl���L*롉b�ط�A�z�90��m
�t�l��A���.��2o3T'�|���7�p^������}z~�c��j�u\��M���z��ck}&����B߅*�8��s�LR��e�L읫��ccaߋ��⋲)�P�@0?����>lW�X��x�6�@x���v����HLa��[�����f9�]������5Ղ=z�٢�����ۄ��mDV�����Q����I0K~���J�[	��Wkt7�D�x1���O��YhJ,�)�]O'�h�y([.V��[�R�O%llE�>�6{��sb�$��ߺ��Ȩ��o>�6}�;��~sA��N}>�w0ϳ��zoeR�9��Yr�.P��nިƋ��+�Ói�z��
�޼���ԇ�����y�D���peYp�F���:s�c9���)A�li�����]hN;�rH9=�X�v��������?!�j�ɂ0��H�s�L;֬�vn2|3߻N{6�p���"rz]�3���O�k�8le��ކ�QJ�'�~���k���B�[��N�^G)J-B���r�ݲ��B�cyO»f��d�HH�;���JF(o>�j�|�^79��)^�U�X�Z��q�o�4b���BA_B��BI��E�%�J�?�1ن�S5��5b}��
^6gM$����y�dѤ�b�/o��D	�E�U2�PÅ0LCZ���hm$�A�Ȭ8�c.%\���-�2� �N��6��_�B��i���ݵ���i���v���έv���nņ��Xժ�V��~d!4�����#D��\��FL�o�m�H�����S�����\l�j���F�UE�)�R�To&�)�ˮ�1���f�s @3�݋x�&X��nl�d�x����tOW�*���W'�T�\+e����}{I)���/���K'6y8��oFi��$�W���X��ԉf��n��������v���%i)��� ��'�Q	�2G�nOw�y�,�ۀfm�FM�E9�zaYL*�8�{?�$]�N��6�!����2��V��(�a����t|5)�������%�l�<�x�i���;���K4,8y7�H��ω/�e/��11AAN���NBU[@�0�WpP�<�I�$s�V�nR����r �@�.�9���;%����ugh�Q�5?�?��:q�{�� �Rt��{/|����@�C�ǺM���P��h��k������<����^%_�Y$rW�b�R]z�w���%}�6X�{�a�u_�]��7$hh�'��r�?��~�t��q��M ��R�J�9$�ɾ2��K_N>�u?^ ��B�1��a)�"�f��g���.b���=��)׽��&L�z��{� 2��j��Un Φ�_Rb��C�n����`t7�O[�D��d����R6���y��ڸ�:i��?�8�l��Ҹ��6|9�_�e�"ݕ���W�M)m�R��9ݟ��3�`��-0���X����ïOY@;w�p^�O�%qi��	U(�}���uLBuk�5"�X��V�������)�p�aQ��%�Ca]�ά	~X���c*H=z�E`<�":)�/��v��֥�E�  �H��.�o�-ͪ��Ra�O����as��J�&���2��a4)����;�$�w_�P_m�&���ck�#�^�uf��~ԝ�+Xnv�O��[K�]Ѧ���E�I�~���)��Ъ ]���O��������TF��z�G��}��j�.�����y��Ġd\�*a��>��a��D9*81�!�L��� �1!i��%��s�-0�\���r�>o"L��G�����9��dnm1���g����A1穛�k���ʿ��o/�G����`b^�+uw|��ӡ%\R�&)�RP�T!v�P`U���o���y+(�� ��;�Ν�a��޲���Z�D	A9��))��$8�<�Hz���7ҪI�u݇��|��oF����I����f ����o�K;kmbN]�Î1�8?��͞�P��'��!���Z��ڑ�	��Y�E=��q�Bo�L�:��k�D����yː$��F��N��fn���Q9�Z���׏$odI��'�c��>�㽚 ?Rȣ�;��У�)����_����z��J�3PoN�x.��p������sKc�Z���If�Ǭ���d�aF�P�B�[_GQ�Y����yFo��T���4����y���7��]C\g�*0t6@�3�p{%WK6���G9'�^����.�<��޾!%\��G���4�z�`X�	�g�}ƃ����>�<��b5Ҵ��:/qt��D����Ξ�C��P.���X;c��	�e�ҘB26��Q"T��MJ(�Y��m�&��)ie�B��'��H�O �e��_P��u��0l�ċ������۷ W�(�[Y���*h�8���f�{޽YW#�_�o~Nm��XHC���S��bm'��o;��2�xIs/�qO�.o\�w<��(*��C}��U.\�&����a5H����v٣��QW��$s��cpD Oa��X0��Y��zϻu�^H��!����:a���������f���|�|����eK�&6��:[���^�י��\���d�w#��SZ%��/���ӴԴ!p7*x*a֝�^�I�k��^u+ק�V��GcM`����|z�u M;fl�󌻙#P��.`$!Q/��f�;�l�үW�kwR~m���~���Z�o�1�����=c���8��ԇ3P�Pc��y(TC��E+=��B���c��+?i[�����V�v��G��-�X�nS�6��\#�N�U���7��� �q���!R�RJ��<C����}��G�qd,���6J��zИt���j�Lm�B��x��T@��̱hC�P}(��9�]�).�C�r�j$�L��"2�mh/��6m}�����'�Y��� n�I{�7���;�UbJ�i���Td�S����SYjQ��f�uA>aq,~��X�BB��Ö�G�4|-�p)!Z��Y��{��!5ϋ����.�w2b⫭�3�G�K����X0��L��=�J��#�� g��e�,ll°
"u���?����'!,��	���$t	�kZ����(�4��k�z�P���5.op���ts�#`�z
��}?0V�9q{������lr�}�6!�n�1`.0��`������Q�MX[E�ۿ��E� |�>2%/N+C ��~&�LK��>��
���v�F)�P��B(����Ԅ\鶭p�:]��|�lrI����Zή�T6�����n���l�N���SԞ>�{����M�Q�QӞ�x$����pHZ<8x>P#o��|7He5A�%c�}mW��6�/e�G�* o|?�D<_�
t�s�3h���m&c(~�LqE~�˙W���#I�<�zd���.)���(��b���5rZf�ڂ�`���3-�Jf�9,�(�,[��1�!P~�����O����L����1�qۘl7�1*��.J�8 Xϓ���4|�KY=�i���o�!��@���]��x����~eV��{�kw|*���ހ�p��dV��IȰ�8}f�Y!{6��K�PX�"G$7�_�߀ò*E�������Z�!�x}#yq-��H"~��1c��J�G*���ԩ`�YT����~�3JD����c�T������% ��wۙ�L��G����S�
e��7���'|�%���,~�����*3VIy,ad���~�O9N�H���Q~�(��P�|��U���;�(�s��6MɜS�~��AD �8�x��IBi��G+�]�9|�w�J*�����ⷴ�4��IOc�n~�0��kr��lPIn��:&�Sx�/����dg�Hw�P�[\�!�)���
��%?{�Jw�޸a�BgA��hY=/Z�P�s�ń��-�~=���c����D�ԏC�4M�JS2֜6�}��������`���t6W�?��ik[-Ì�~
�Q�&E^���61�$t�z^t�'���N/����YZ��`������9[��$,;��໛pA,����K<���z�#-I_�Tҹr�� ĭ��h� �q/d�er8p�;��ʴ��%��Wa�Z�~���P�j9ʆ�f��-�E�<��F�va찹��)���@$��a,a&u�~r��j�	h�%�]�����@�$��QW&т��롃.�_�{��4MS��'�C����P�6�P[�oP�sY�1��8_j�!NT���^|����;���0]����iς/o��Y�#�$'��\P�"<[��~ w�~p�7Ӕ���Z���jh��O.���`�|&(���PR�2��+kh�%m�w2�gj�>�|��t�`�n����b��>��A(ʕ
be�B�A3�X��Ec�o��+C���������(sz�˓-��՟��0�Cp���)"(G�׈���4�����@{�`�����W"��V����o�"�%�e����P��}�
��G]��d�^��>�0�x���lk�1����Y��϶�8�@�?�w�H��T�R�܂d���ų9Dv)%:6���`:ف�,yp�8�h�u���4�}rĊ���0�S��}�ߖ}���Σ����m[��O�y��h�.���M	�0���#IxA�Lx!3.�-e�U�6uyB�%v΀��3/M�60��zF�����}�J��¦�G/��c&굹�\t��&���z�L7j�u�m_J����rT���Ws*���Cgw��a��� Z��?����/�$�ǂA}(����p��������;�������Ae��!��<р�n橶L�o���T�h��[���z�S2�,�&D�#�-�;<�	}x��Ȏ2�^�
(��/_�B�`�K�O3�O;����oH��r��|5���ѿ$d�ƻ�R'HД�X�˙�1��Gܝ'������}x_ʤn���-�pt�.�M��r�Npm�����i�p���)9R�3��x4v���h ����.��u8�SV0f<��Z�G�X|{]`ZȠ�R��l�ws2�9��;ng�p�h����;t!���赙{�����[Q�+�������#P'E3]}�8�8�]�t��B�|�:�[���`b��E�#���t�^k�f���dHߧT��)�궏}5���_{�9�@�@"�6�c��d�i�fϓ���Vw�3	"�&4${U��g�>_�/^�,}�zlnzLn����PT�>�P����
��v�����. L���^���7i��ʬ�E���U���v�^�-�^G9��佡��zT�?�ۊ���r�˵��8�D��:��&���y-��>�ԍ��5�������`G��z	Ί�f�a]:z>�k��4�
^j'�Ҕ�_j��W�k���0z{NP����F�Ҵ]�~�GNeJ�,פ^1�`}��,]�h�ilعT�³X�K���5,�WѢ�����C���2;�V�����M̨��/��IF77MW�4:&+�D�BXo��|eŚW������{���Y̽�_��6������(�ƪ:���l�}A�蜹��"�w��G�ö��(o�q���ø��J�e;���g�����%9�E*鑋<��ؿ��������R��v(����6D���A�>M]?_F\�ǁ[��He|��6��J�M�,G3=Iύ�ݴ��;�<�Hbo�}����MGEe��*:!a�>�n��1���Ѓ;�ŃJ՘��>ؖA��\�c��u��'�&C�M��qVtY����hx'D�>!�6�}&���J��$Ю9�U6����z���'E�u���X&��Re�}����	k�����j�O�B
ѩ���v�6a@�O,�g,?a��g��i窩�/�
��|BSL(�:��"���<%*)�u�z���0Ë��͋�q�
��b�1j���bg���9`����{�e���>�N^\�M�o]��c��_x���.d'L�N�q@�Uo��RL�(6������64	 |֒~�k>C(��0Z�j��Ko��+&�=�Y<��t�8#���i��?�\M�h��b~�./��'��4]��a�F�7��Ry���>)�d0�9�ǆ��� 6S�O��WpQ�;��#��f
�D$*�V��-W+Q*�_F��&�u$��/����[�K�❝��m�߮m��a�5��i��H�����K8�K`��S6��~s�����0g�	u姣8��[(,b�9�ۍ�����h�}��B����w
!*� ��yg�eD �8L���px��0�6VU�A������%���y{������HU2�<���?X|�
��#�T�d}�\<n����}\��8Y���-�;@�T��+O`������WƟj�a�3��@�f�Ӻ%4�����Z��C�{�>�'J��o,���ZO5����aI^o���J���j�]�U҃��_7]������1/���K���T5��4����09,�q����<lǕj�%:���-�;_��� n=O��L���t~�:���e	��x���6�~�(3�'GE��n�k�I�p��_5RP��H�@l)a��{�!�Z��]l�y^��?�6�5���.L$�i��:<YX�}��=k:Xu����2Ǖ���.�4��o*��b�Ų�L7�f�Z[ʸ	�����]'kў��)�6�2 `a���ν%E���O��*�C�.:��'g��{�������,���Q(�7�8�Y�V�����ѻ<�[�0�xX1W1n�BQ�i�{��ݼ�;�N��1���3�jن������c�s�`��' �l��_픐\���TZ�8�W����tr@�T���ےYM^蝗��������(|6ٻ~IH��,H��e������^���¯{�x��Vg��e���Kw ��VO̓�JV�\n�D�A�4��������ڴ���:�*�E����>�*�>�xR$�f��m��E�B��}�<��Nr��ʾ����`0��5�\�F�f.����S�:P|�?��Y�Y�����K�Y� �6*mY�Vry����1��N�|T�2ܮ�u�d�9��:�sՂ|��ec���6H�p-fBۅ`���1>FW��t�����.�0���10n8��~xtY�6u>TխA� �� PΗ�r�v�'�Ad�ү��c>�������箵�,X�6�B����H�VQ��=7X�<�C>��͒'����6l�S�+�M�B=Ѭ�o��,N���B�PT�+���.OrG�D��=��p�2\gp��t�xmAe����d������4.�u���Z��Sht�r���o�3Z�Y�"�_Q+1dU��*#3척�P����h��߸�/���oo2kc��Åb�:�BN|<}���|J�~����:d!�0}�������
��/2������-���W����I�Ͽ&+�m�y���h�#pL��@��f4�3�:e�fg��o�%O�q(�%��Lz,_�5�@K�ɴ�Ws��9�H���[Y��4 ����RS��';"���a�#���05��C�z����K�12��׌���;�/AI�q}�<?T���Y���Sp��9#��F��*To(; ��<Q�Y��n�D�\�G},ڳ��MU#�5rFM���<���RR@�%��,o�q�j����)�a�<����Erw���ne����S/�;\��n��r��=x�*$8L_,��sI������1���s-c]�o����ᡸ�-A�\*%r��?[>��a�s̫p��4v"0�����g�r�8S� ��=�7+iD~���F�6=و��$����Y0MC�:m��WX��IjEm�<h�H7:\�t90ͺ��+�h��H2�C�#�)>�E�{�/�qŀh0�Ԝ�nҰ}�R�b�\����:�|�$��G�����:�G�g)΀��2j�P�|��ߚ?�R��;��k���S�h�vc#��I��*�7�*��2�}��)���k~���sv��a�N46�t� ���u����c��0M?g��6] �}dW�S�vf�{�O��.͚�2S�ni��7�F���.�	W� r̸��V�@�0��R��Yȴ��Z:�W?��.Y�R־�)m`�\��U�n0��|`��J��9	�9��m�J�I@L�?���\)�FL��i�jz ����ko������N�4���TӚɶ�jvEfH�_(�/��ݭ����D*t_F��ڍ��,D���	�ٚw�/hn11�6�(��N��<ccz:�a�������n���G'���01vO-_�V.���?9$}���})3�	����K3l�r���b��)�Cd�J�^_��C�^"���6�l1�m9a�I-C����Ē2( l�f#���`"���,�f��-�o/��M��m�@�U^,�;y��?���d�<�_ݻ#�5*�F}����H���:9�m���'y�tK��PD�����P!(��*��v�S��%zG��8��[��;*�!����bUkf7�d�ܹ.։/���"`�_���%�2��-����˅�=~.yC>�\�����\�'.���=���V���`YU�w����5	�@�uC�skn�3\�Ff�-�B|��s�&y/F�䒻�8�I��h�2��h���q�#�0�3�$l�x#S�fÝ�p��sP`�D�#v*�eR���!)��q��� ��2�Ɵ�^9d'�I����� ���͢n��b������#������[���t�J�Mn�6�n�����*��+c�ﱴ{����QT
�UK�=Qt�NP埈�2'"A
۳��f����.�7�\YE
��x�s
$���"U��^�E
.�xwBe����jP�k���)�U�e���}0�����D��
�ȭHT�>�u������D�ן��l󱿭.z\�\��S�mwy��b��$���R.��9�z��|��;�7��'�>n�b�!ocs�<J��N�
�iw���~8Z�7�=��h���E�(H�g����k�� tg� ��]/#�{�-�$͘�����{0Z��t�j��#2`'���[ok,�А(5�� �M��Ot���Z� �]��N}���C�ȧN��!4]��k4��	����vy�[㕁�)�6՞.�oE�Z�Mt�����P�Rv/�%̹*�u�)yC��'+��'�E��o@υ��X��Q�P�
Z���,�?��?�-y�|�xk������>��Fr��<X)��P�O	 �����h�%o�>�%���L���n�mQ�[��;�%`{���"e Kl��Ϳ~y�L���<Ĵ�3c�pF-3���(K\}D�)��ɷxt��g��"ah�W>�����s>hr	U��OARx2�4�&�^�����5�&	���bW�G6k�i��c�ɲ׊�U�8\X2q��ǔH �-+|)�-E�#��T��B�2�F-<�N+tL�Kr��;ʻ��N��v���fʽ(e�B���>���jb�	���1���(�����x��yէ�^N7��Q�F� �bL/��'5�ȒYc_څ���K
�5畄$u�nbP�ڕ;��"C�U݋���)Rʭ
���F]���<!#X}��K�D���3>��;�^q� Ƞ����B��q�n����aȝN��qdb:����)ϰ>)�ݲp�@�~2�ٸA�Hu�"���n:��4��������&�>�0Ý�k�pEK]��]b�5���N�dFޛ���L$���0�:����5���۹o'7%W��K��4��A4gyY�E�Ώ;N�:��f�5p����2A����M
y�gt�����6��1��Q7��>��Q��r\���^F�/�őH��b��Sr���������TG4a8���1V�S��U�o��J��Ⱦ�R�5�w^���>�/�t����p֩����+�w�
N����[˴L͗����-A����Q��R�I �%��N�wVրXy �
?��L�%8��Oi� k����_�����r�T:�0iC��u���F�Ӫ%����'ԉD����z�E�d�"|�!D�6���2�}Zc�S޵9�n����mh�gHΪ�qs�6�G~��QCC�����0s;X@�W�7��+�m���h�A�Zj�L٬H�9����
-k��kM����'�Xs%�0��.
2,je���Ʀ��7.�麧5��ؐR�]Z�$k>���G	m�j��q�_#�UF�Ԣ8״�"1u3)�7�i�\C���o�u�tNkH^�q^���S/��"4%�Ӏ��m��d����G$)�������5Y�p�)���ž���^'䩪��U�u���<~�N�|�A���b��?q8%.#k�b�2�$O�1�<�!���C��|aڡ.eo�m��m�;ᷘ�)���e���+����L�����g(�2�Y�6��`]<��sZ��"�ӂ&-���C�-́eua^��{K��f�z� ���҈E�3h�6�R�2�R̔~������ 2�����a�(�x�b&xl�v~M�c4���1���E�X�g� ��� b���l}�PP3)����:��]dZ 5��@�[H�\H�G9�U-���jÝsI��5*6X�L�x?��3�ni��<��X�G���㖮jn��f�(�܎*� �W;`�����T�]����%��*�����ǹ ��0�i�$� �;k�� 0-���uHf�/n����A�"��y�$ЭOF�5�����+��[�����s�"K��ү��b�."�0׳\�
��+��1��~U�f�k�䜀��4��=J���� ��lF���v"%`�6���&�9��Pl(.~4��[A�1|�S�����~�/��|�7�7�A��?{cY�~ε݅`�!zC�!4�2
*�G%�����-������{�*�Ὺ�H3��fǤ���/�u�rؒ�X��Z���0�R_d>òZ����i�JXb$- �r��Aeĵ1�/�S�y`��a����;L��$��K!&��x�zm�I�o#>X �.�U����J�@e/M�c�7\M�ї�%?>~U|Fx'2C�L���G��Z�F`����t�����z��c��_?���������H��p�,�fK�g��X5��p���o��-;�1÷�H&R]$���I<��lVn�JAJ��N|޷�,��J�D�N���5��>5��������xu!� ��Yȧ~8��<ξ]������ϳ�Z�6���{+�ܬ�����	ƃkyzQ�e���m��?z��A����ѝ`�� ^� �юXё7;0�س���
��kݽ$�;����Ш�ȓ��z*�ߴS���F�\|L���e����PPe>2�p��71�d.FP
���
F�c�!+���lܘ��C�+/�����{�<�����I�~�,��Z��m�ڹ���S_w�D�KkTu.�7�C�<��s��1����}�Aߓ"�*���>�X������u�����x�5�n=���d~0[Ԑ`�x4)�J���.vIŷ�=L=i�T��y�3eP��(y섖��������.��m��(�cf��X|�i}�܀��e���QD�@/�1Ĉ���Ӷ��e�z,�����Ҝ�(`٣|�SPv#�i�p(�>�-?b��MA�u�L�u�>��*��#��}�2���<�նG&w��S^��&��Y�B��d@��`w^��|�7�%7��/��U�s�L�8���	�9�i��mi�k^��P18�,B������Wa����}�h:���b�\qǰ�pɂ<���ެ����@�n�;���v���`�WUV¾���DTr��U'����T�����(D��0�
�G��z�*(u`k9�V��N�0zt�̯\Kc�:(3vKZ	ذq�X%�.�q��0v�L�C�լ61-��70�T#`0����o�%l�dU�!����2��OϽ�/qO�'Em���)�0k�+B����yS/&�z�3���H�
&���X�0��
��8��M�@�����V�:�X��>_�I1.��C��z��@J*.+䲞�9Ǫ`AƠY�w}�,�Rn�r:n�Ks�N���7�"�<��̥>r����7ou������!��=����Մs�gzI���s�"U)ؑ�T��'|�,RO��e�g���
���sJ
�'r:S���y(�k!����6��I${c^� �� Dd���}�3��32�4
7Ao��8���C���2�M�?a��i^T��ȼ�Dr&o a����h�}����F��I�XQ:1����Ua�^��@��6�ȥH!�osy�"�����Ԫ�+gK}xβ7�RF��"��;�,'e�48x48���)�v�dqǊ����*m'e�MB����ߠ;I��7<x�IS�σ�Շ��̻�Z�İ!8���מ��N�����n�L7r��j�:���'B�S�}�&�zݍdTV����7�ծj�8��{�|`�j ԼX\�R�v軻����\�k��<�v'��}}U��S6H �ر����k�?G�F��f�	%.r:���o��ʫO���#�S!�3�a0A�J_x��W�t���g%1�Z��j���-6�-Q�$z��e�=%��R𹰳��$,q,�f:��?��=�E~�_s��j���)�
���̕-]�%���W��<].�����x�� �$�5cs�')Υ�94���,���f9�e�'���n��Tj畓 ,��ʫ����,S,QȘ���X�a��!}@�/� A�Rv��f�%t՘	c��o� {��$��Wcĉ�q�A������
I���k�T�3���t�x���m`�!��׋������Z��OH��WL&[��6��
�Բ��u�
�au�_����^���#m�,���,C6H]
�!K4�T��o�0	�n����,L-���nLA��k1��c}\"��g��C�4�!��&������#]�y�9Bbp�I�wmf̭���nP��9��%��7��*�JP#�g Ds���������ڐ��c���JsȎ'´R����M&(�P`�!�MݱK��D��128�b�ݚI7�D�����ΰ�A;v�)��)4�V�&�[(��6R9̐�"�v��"�5����?�m �{֔�.FF*^{��a�KkWp��$^q�h�if���"I�z0"��R&%���Y�)��\ݲ�B�W�l	���<7gtU�*��D�U�˞������ad�:����K����^��CA�u�t���o'0��*u{�
N���|t�Ҏ"d��T&�vz%�û/��O�8�-g�9���}��mkT����Įv�g^���d_n��˗���ug04?|_u���܀ov��@��:׽E��?�OO/�Ӵ�6�����J�n�C���Uߛ���8	
�sV�d|� �5�b̢�B�fP�P�ix�W�73_�C���G����'�uɒi�J����/IC�B_l���&��_C�f`
�2���@O��_�bE�=�-��/l�j���]���w��ty(��A�,�W�I�q��_X������N���������#��i��ґ�̱����v�}*�}�ю��qP��ColG�b��X�ʎL�@V���Q��d+π�l�m�ћ������9"m��H�'��vP�'Z<�+W&8�h 7tE\��]#��n-"a��[�1�'�-�ce�Fh�F�I��L�vn_^���>��X{��6s
�Y4�����]^���{�÷p�|���Ǩ��f�QEl�z����HH�\�޸��U$ʄ�t���)%Bei�
TcD;Z�M�G$�l2?x9��4�6f�Z~��7��SÅ#�³��v�J���nE��������/&��  �Xo#�� Z�����޴�]N4P�
�����Ï-�Km[���)��U�0ִV���~����TF� ����4M6y]ېf2N<�U0���L��P���^AtZ�d��A��p'ӵ�蔮Rť!��p{,�����l�z~Q�r� ����������D7�:�=����i�Q#���N.2h+��1�V)��QK�������5�I#�c�oէ,!��Vj����`�f��dZR��d_nd�]�g?iH*�wF�{4�w���,6�f?���dF�k���&���ay�{]Nf�ꔽ���ֵm��ʰ����^H�8��>~5W�B��c0��ƪ2Sŕ�{���H]�̊3�G_�4�
�ln�V���O��V���2k��M��ɏ�h��D���6jR�S����eTB�a�]I&������2��mi�kvv�ŀ�u��"����<RhmN�����I�I��MF��Zw�1)\k�`ĸ�	h5�XE�EW�]�1ɕ�M��t��Ǣ�/	��8ƟJ��+AM ��TБz��XZ�:�z�]��kmX	w�N���G`�W>t��B��(����}��R&xぉ9ƨ����<�����ʤ
�%�2n��9e�_�.5	k'|����@oX�X���߯q9�8Lw����Jc���fZ᪀�^�+C��;N���f�@��c+�Ɇ�l�=���Z�9 ���}����7�lq�����CZ�L�&u�"�G�4�=Dܪ���W#0)�X q�\-!)�1�K�.������a����Geⓖ��E8Cr��\
g?!�˫��c2�'��7q��Ҍ��C�N#'}1DxU��gۚ��K-B�RxN0��pP�z���\8�yȃҧ(�K��j���
�z�������Q*�C�C.}�z�ե�8���������1%�s���eM��j���qWbmy����_��m��^�6]Ν��@��F�aB�-))ə�l!�*�$0���!����ݸP��LK^�`��k��Z�1��<�r�����m5F�.nglFݍ��z�G����J�`d
������iR��bvI�_��:1d�&��!e'��NH���3��QJ��{P"V*[���M�w��	Ki�2fXj�=�K�2d΢��dy�pG���IF�Zf�n����d=�p1|3�bn�i�ĵ��k�T�_@�x�����P���y��
�f�LQ�~7᧭����X��5�r�!��P�nC��5QW��;���\Qk���eQ�QK�󉞙q�����|B`&��5�_�GC�)s�w�����(��Ġ�o"otF�\J�3X�1�^^8SLwH�<8�,��1L��`0�:v�7Wz럼g���6�̮�:��6������6��Zl9�1���㎹���|�:���L�9%�:�4̸H��Q�w��:�[���u���ۏ��n�Ni��g��(�UxRh�!�8W��F��&Y�0Ⱶm�:6
F�6�$��Mu`%h���Q���e�c�'�����t(�ԣ�����R{�I�r_��@�ji\��E�{+�ϑ��]�ۙQn���9���Tk�l�M_fHM��S�j�	.������eq��:&z�u���fL��S"�v{h��Cf��S3L����A��g;�܌�������lxJw}C�$���	@��8�~\??ԸB��]�D��ݰ&]c��j<Z+��q�u����=M+3��_ƪ���՜������d�zC��ʃj+6d()P^}��_Hjo�j|�~������xS\�G��e<���i>)�[��>�f���Q}o���L@��}�,a���b *�z����ld��?�n@�����>��t��,��e�A��+��p^@�A*T���c��CE8 J���~�I��Ү�����x�3[w��	�Կlݼ����/f-�J����B�u���`�?�G�b�[y���^���U�9u���$Ώ����@��߁�&�&L*Q>�<G\���]�T���d��2|�bDCOf~w�hKEQXb5�ݵ8�m����%�C�U��(���RX�%�U��g�LEX`�χG�'#(k���Zv��B��f����@F�X��!,��ɵwKD0�p8k�#̚�u��?���'�2c��v�.��LQ�c���ḯ�+�U[�Q��{�]>n%��Ŕ��g�>���{���Y�$���Be~+�j�Q�=�5ۈ]��`�s�Ĉ� V�Z�w����V�Δ^���k:�!a�2�9�!��^�/^��T�� ;�CcEA��6�N�b�5Ŧ2ytp�+P�4O�V�:�q�K���笫R~�Y�RHC�y��vI&Qe��Nv]���@l��Ѳo���r=:�^�O�:v��jq�K�a�9`��?�i�A���L6{k�2r��Ea����}��PU�<� Mӣq���}ӽ�mR~�h�bɲ�9�/AT����]��]<������ɩ���G �nrY^~
>Z.me�DM	|����0Y��l"tçH@�����]���	O��wջ����׮wK������y���`"�:nf�ڣb=�!2��;��4�F0�\�����[���0�f�_7�G��h=�9 q5�M�9~�A��H�-�b��ѭ�(���ޭNV��yS&�s#q�h��Ȟ���@�*T��c�D����4M�%����Eoܱ�\e��	�.�IJ{�4[/a�vL�Q��:�e[�k�}b@��n���B�����lA)5%I�xT��8>��d�go���P��=�#���^�*��MkŦn}oC���y˰!�Py̌�E��КV5�;&r��
���vBl��F�W"����O}d��u[Wظ�ؐ~O�����ݷ�;4���AQ�iM�^�YkO��(ȕ���|]��Ie�?Ƹv�S_n�qB��N��EZ��겓��q񓮶*�+��5�s.K dM���~-�
`QAv��a�:�&f�{1G���*��q�RfO5w�o~��H�ۤ�KΙ�+��X���s>�����N�]%��K".��F�}�j����x@��@�w�?|��0:0z[̤b��U�dO>GPi�?l�����T��,���^.a�g���ք�����Aܳ��g�^D,0��z~f)IƩ��9��ޑ��K�U�R��{��
�[���]�<_��ɌH	�K��!)���X~M3����d�Y`d!�<�w����O�L?���lP%k��(���ض��[^b��R�#q�L�>��]��\S"��O�Q��$��D�|�68&�=�������'R���I3��7%7"���`�^��g����+m�kS��"�݌�}�oA��X�>W�M�<�4������À��\��:�WnhxW �Rhe����&�\��4�9����G�{�̶'��k�9�8�[[�_���S�\�;Q9�/�1�P�Ҹ�Q0�T���"?o���G��wh@��<D+�Ч���jLN(�W#G^��O���5���;��U�U���Th�	��'@���mٜ)���I �� ��	��H��	�^���D����������h�1���{~��~�μ�����N�J%� ~����M� ���L�`�)�8��p3�9��W����ɉႾ�~�Ҭ�{r��ʊ�otG1��e�F�а�I$7)�e]��:��L�7O�sBk��zj���(�?��g��L ���;��}mS�h
r1ѫ%N�]i��5�הk}�䜻�h먤�
���%����b3b�d5z��WV��=��?b��� o(���ӃF�x2�,1
-���8D5D�A��=��F���l�������I\�jǫ;�=~������$�t���e�|�����\5@����?��YS��d�m���'�X4!����/{����ث�׬��@��[Ŕ0����I��0	t$��'$������*$�ެ�ʇ�u`ޖpCHB�$2	��m~	+�)�C:��jGt<���&��̃�/��%����ٷ�aD_�2� i��Fb���ň����2��B���`�,u�ӻ��Qc���:�߹��RQ�R^�k�D?��d�|b��UM/�\#5��@V��]�x懍9-jk�y��.@�h�j!�N>?�G+0!�B�xw�?6+��{�I
E=P�c� \48?�-�}fj�=�I�:A�_�' ��ܖ2�5ڒ��4>I[7�ۂ�r�Gt���H(��U�udb����X���8�w]y7�o���Dך�������=|}�:����'!�/�nYL�� �����*@D~�z�au�(rm�����9+q�6��1���j��(��"%|bl` �bA>V�N3)o�sJG�(�7jJ����i�6����̡����1�~���ӱ?F�� Z���E]=N�R���� Ǒ�PV:"����HN��ҏ8m�4�D2��j�>�,�0�n@̶�]$�{�4���<�Ϊ[�x|�${^�x��:�����L�NAU�Ŧ^�9�m.Uv����<F�������g�����O��!���ʦ,pQE�n�0<I����O��g�~W�7�^*�1F�)��7�ȝ�E{�y�!�� ;�ՉЪa=@#��4��Fѻ���3�����d��R�.f,����JKtd���mq,w�_�?���즂�_��������IKnѕ��
�R4)�>�5��W���v��$vkPm�sJ���J
-�\cfX����7eS1 ��`�H3o%z̶ӽr�hz_j�m�H$��o;T�X�kP��*�߈t��/�k�l) k�r9O����ً�T�
����R�tRa.�I�P�e��������ǖ�l�˓]���n>m=9�J䊣��&cUВ87��f*��;��A����*���7����~c�n�l��i��d���B�4D�����M���5v�u_CmjD���Ca�WG�EէHqm~+���>.���![�Igj�)� &�dᅔ�&f�9&07*�6��*��� ;%V6��F5b3f	Ɩ��/����@�	�����P�R�������
�z�w�d�8��e�K��7�}iX.��l7.O�tC6���ϳg��I �s�)�<QߥA	&��c`���� ���	�v҅DX��Z	p��J��D��0�Ϡ������l�N'�n "���-K �����x�� �*��[����¿�ț�8�+�ի}ц�����׺]S4����E�&���ӯ�.X��6�4����CA� ��4����3C@$���Ԕ ޴0z9���-�(F���Q`�D��f�N�o�R[ԍS�>�T���Ȧ�8\B���.3� �M�!UF��n���?����:]�AV�Ί@=��C�����h|�6^%%T����D�'����p�c,˸\�x���z�L�(����K�v�M����l�Y2�ר�W�ķ���]M(�ŮQ�+q8��]��ҽ��D,� R�*t^hMJާ�P<ae�i�ˀԑ(��v�[剏^Y�
��(�
��un���Q�=�%�U�G'�2����1�2��*�7���"P����ã�@SB���ο�=�9ȃz���	~ɭ�G�����uC���Q����+N��*���~��V�N*m��������f>ͱ�^����F�[@f��1���b���H|]�h����5�t�^k�"��8���m�c�/#*��2���=�z��KN��W��tY�1ƣV��l!�+���I��ے�F/k���]sDP����3��u���d�5��YuY���"M'q*FCH�T��INdͼۣ�O�C �-�"�;�fq������+� �j'pZ�چ)% a����>���j����/��`Rd��*Yt\j �V�ff�B�V�k�s��=M'@FD���5��l`o�fOcLnN�va�P;� �57��Z���
Uc����vr\Q�H�����bf'������Mu�Htk�z�1ź��j��;��nK�i��"�R�ﭶ�Ys�.߿���E8��qxw��҉�!���of��eF�Ӹ���o��9����r܆	(�a��l���		w��=D
�U���.Ҕ�ct�o|��"�/rϬ��{DfM��i�5	�C!%{�aee��~��&7�}�n��"�O(��j�UG�6�� ��O~�-�kqy��8�|�y������2�e��Ǟ]�a
��@8���ӡ� i�s��VFp!"o|U�MY�'0���%��2H������Rh��ё�}�!j�.ɇ�|#�}M���KO-E�(Ҋ~i����/7t9H8&�4E0�tG^8՚�+$��20$�̏�*��|MY�?��*o`.��M���EY!I�؊<_��Ϟ��"�nn>�[�CdmJ̆?�-\�ߦ���b3%�ihe�;�e�Cȣ�wV�呾��C�ⰱ���"H>蚎2Vƃضkv�±!�rI���ߐ��:�bc�dN��xo�9���{Y�Vy�l��a����Fq����:G*�C�E��r�t|�����CL�� I8�)�����1U'-�q��,���D�/6�׶5����I#nZ�(@���O���t���
�G�.i��q�}TH�b�߁ۤ�ݠT5@�G�M�83�y�t+�~Q��T��G���w�����d_~�7%N�>��s�[a�>QvB��򽡷n��BD��4#��4Q]��0q�ɘ	ޥ�m��+B0۰�d �w���#�f�E��dS܁`J`n�\̤Xar��9u��L��LR�Tk�v�G�"1t$���$��,���^���].���!>=��kB́����z���o2���`)f!"ug��N̕�Ft}
��#p�;5�#���dzw�9;��%D��ǧ;�!�Sah������P]�뮣n�9��y�מ�p"�t���e���w�Yw�~�R@��zȸ�v�\\/o�ŋ������(��y4�����
��à�+yN�S!֤�Ȇ41y�P��$S���l��@�@.q9�(mZ.�(ވu�v�IKz�8?���M����]~VN���L�}���ܲ���@�i�;<�g��$�����O�D�J�G�E���5e�!��
~ߏ���v��?�$��f��sa�ck�����+����j2v���bl��w��9&��qZ'@�X�X7��}��~B�����>��s�l�iTp	yB��x���T!Q
d*���e�$�~*L^��ng$������5��#��o�&�b����}d�0{�f<��,�K}r����ދ+;��{�Mt�)��i�}���_��Y(� 2�{8�ݵyT6�������1}�$mb,����0�Ӷ�\.f3��!�7�� ����Ko�Rz�l��9�J��l�#�˭�~�+)��ӞeC�Y��$���k�09��x|�SP>u(j'O&��xc�cI��s}VſW�/r���U��Y�ԅ�q�p%����Y$������v��j|�D)���i�:��8:��'�X����c5�Pl>�'���f,��3��9$7FT5�F����H���2�+��=hU���t;��P�����޼� I�cd�,mOT���Y�T��%� ¦F�>{��p����T����n&3;�u�`Fq�熷��[����s���f�e��{舷fq��&)�(6��;� �|L�>eu��DG��|�C���v�{���w�"��e_��ʑ�y+U�aw9��`}7����{J�ұ���	qK�޼m'���"�+����y��(Fj�E���iq�\1yW��$��VΕ-pXmES��";��ִ��x�L+]➊�҈�]%/�Λ�˱<6��g�A#6i0��'�j�/�p8���D.��s�^X��GN�\q�.�fb���6ؚ��N���'����φ���ĲsF��2�\{�^6xu%�n�Ë?�'�D��k-�9õ��6ր���2 ?��*M��{������yb�� d���{n}�Ʀf���,p�}F�S���G�S�>��$�?���m�W�Z���7
a������8���a~:p�X��VOӖ��>�m�"���HJ��u�WNO4�z�bSb{r�A��IÌ�]H���s)Ϳ� ]�O7�G���Vq�)��=��1�N�Z�9������;}~�n�6��M?uj_vJ�[>sZE�Ikz���B�z�%���<ukD�>����%��Q�R<�y�tm����.���3��n���#��J@���Ջ����yW_S $ݣ��,�q��p�6|i�����B>*G�e�~�`:�2.�=�+��Yڇ��
]����Te@1�����$�K�i�9̚JQ$<A��īm�\�1Ƕ'׏u���M����4�C�I�����ǯr��\��Ɛ�#������u(5��l'[��$cT��B�P�XB��\�%�z�6b��M�wl��y�;6N��p�=P|��vwijc(���+�Ǧ�*(<�b���y;{7^���"���v�����_��l�`����Pfr_,�`B�V�Q��bIZա���>F�N�#n����{�Xn��~c�#
�����Xh����XF?�]C�vCN�)�|�[�H��c�Y����\B���e/¶!Q�Z��K��h�0��0����w�kC����*05X�����U��c]�'� )Q��v�g*t�n�Z�!<�9a�$��oep��qEJ݉4�.E�΃�ϴq!�����j�e0�v`Yޝ�%�,}��޲Q�"̆���,^S��S[��jX#�l���w{�b������΃�z�DY
���iqVd5�t��㹟T���?�0��u��W�IHF�f�p���w���d@�����> �%�-�;L�!<��z(ρ�滚��U~�)�-����b[	1���%�n[�)%W%�K���?���Y���)�n�'G��JG*��+�]$8���p�i�~s�#]��ꕛm��DC[��#D��h�[�L�S~�W��ǠE�����2�UjSG�d���B�$6D&�mY��(Xd���0�w��Hs�����)����:|ɉ���nC1�m��^ZU���&-s�G���]��ro;�*��R�z�Ѥ���kY@|�r���v�=�a�v�a��]P�Mf���]5e�Rwsx�&*�3B�~`��+S�Ę"C��:.���A�k�L��K�B�'q������{/>;l0c�v �le����)I}����k���k�s�,�K�716u$�/���xuե��Zj
�mt�Ym1�+�rEY� "w����F)eW�׍���Ş@l��}h��'�c�R�q5k�g����nvh��c����M^��f�eȧ�&�k�Uޒ}]"+&�1WQG����H��N�p���9�PuR 	{ ��g�}�QT�o"��?q�T��I�d�(j~��C��>9v�7/�߆��2H�s�BlQh��D�X��ܰ������|K%g�N�ru�+��n�t4/@r@Y��4~\���?�q�K�^,�LNe{b�-^�EĘ�x=@A��:A7!�q5�m҃���QQ"�k�:�%&PV���X�`�A 83Nu��_z]��C�t���uq�?������������i���4�۵��9�h�W��y�'�V�H��� ���ڀ6�x�ƺd��R�剪�=�a={'�$�3�-|�%I�C�-	�d� �/����@x��_��o8	R4t��p�d����V&�-�t���O:�U';��!�c��{���\�>�!R�a�
 ��E����5��½�i�BVȒ+�dN�f��z�_3��g��)�3|�c��*�'os�?�ܟ��9W4}�6�y%+`Gu��{r���i�����������>(�Ymj�Gm$���PM�^����hdt�����V[ߧ��(P/5�m��.u`���]�D�$��)�\��J�*ۜƣq�Aм)ˤ��/�v�-Y�ɣ}��!#b�����&�G_���$��o��u�oUlZ��������+�7n�^U�bĝqVM��cTQ�G�d+��Dd?k@��>ᐄ{f�n����o$�P�K����|��B�^n�Ɯ�?z���� (��.�1�?0�(s��o�j��Cla�華v���I�OZ�(f�_�cc��2��Em��ǩ�D���>.@z�  r�=�W�6��o9(�`��<5p��KcL�p#��#�-��h"�˱��<4VMZ%���w3_���6�w��+��\����{��͈�ϛ��/d�W'��9���o���iJ�+W�'��ԅ?�oOsL�kHJA`4��z{�;��r��Qy�+\��ל��	|B8jd�t-Y&�������}�躁Fw���c����M��"v ����6��:<��+������h�,���y4��C�˶gZu�������d�\�Qf���B�{TL�!�%�Lh#��"Lf��`�U{��eI����������I�AD�����9�tR�z!y	�n�4kzj����&�Y�5-"џ�����ox���H�Nd������l=���o@�0��2Q��A,�]�Z��t�D��|Q�դ$6B��.>��#�Ӫ�J��O�5V�I(q�[y����̚�}Ҍ�A<�.a�2�7qj���ץ�(�u�^��teR���ځ�J'��g��A2Hxԗ��ɤK�j��nXD��r���`,���vP�L��Je���,9�ʌd:���-Ƙ��Tm� ^������9-���dǾNt/ˇ��Y�E�ɢx%~5Uӫ6)�-'�^��]P"�"m����9a��NH�3�\��R�l�Q�Q^޶ZZ���L����W.B��G���|UG6fCDs+\y�{s�w��KW7d>4� C��u�o��~j�>ց2dl>�}��%R|D�'[,���r�,0�Ol��/F{J��R�t8I
���,�ӭ������9է��D��1�j����fP��듍f1��;RM�`�Ğ�<Q�Igߔ':S�Ą�boV�@�L,)�I�ǒʌ�F�(��˯*+�+؏*�˶ͫ��E��MQ��h��f�WW����D���3�ߌt��U�:'y{3��p�X+b�BS�K�*��`͑�*!����c�P��@M逭����ƞ���V��s��������YT�w�ﺹ�E8	��+fϸ%ӪY`Ֆ�0)��i�oX�9�7��d��/z�x��-;�T'r���I���͝}�ù��eG�	�@Y��3�x����6�<�����9R%���o3�F�L̎/$��{��Ł)��6M�e���9�*�r$��3�Y���]ݞb-�i��3C�6�_���AY"aϳ��q���3���_ƟɈ������I�<�l�4�aA,K�>�B�k�lL����wPꔻ#d�r&�-PjڵAU���Ѧ�m�����pT�fhh������)�bn�k6�Py�d�����_�ø���5��hO���y[i�r�b�;�KzX�ԲOf��1���X]�vz)T��Λ�MB%��15-�lu4B8EЖ�aX`�$��VF��\�>?����n����?�r1"Й{�X6���:��D��կ5vk|�}Տpsc�}���)��/H����n9��A����#�Ø��b���e�`H�jC>�(���=������NVOS�R��g�0� \W|5�d�_�o���p��J����yv��a87G_�kV�7×�������G����Q�$P�QW��ʮ�H�ۢy�7�^��`�!gg?G�ɋ0h���Į㊔����-K�b,�ސ��5��V�Ce�X�.�(��_
'�,TH��IC��1Ve<��\f�O
v���P'��g�a#����B�R��v��k-� A �f�g�|��Ƙ��%��V1M���N�si�V���Ytb)�lp"���q%�'��;�^v�`��V��:�0�����)�j�RU�����AӶx��f���ri���eh�|_���WYhѹ2`�/>�(E�����V�zi�'�t2�2��J!������
e�h���s䑒�k˽K����U/���#_2�О��f�Q���>�&ɟ�׶w���ص#Y�p������3����#/�RP���7�Wf��p�a���	�a)��$�ƨއ ��rܒd8�rվ��I�iV�I�-�\�g�k�%��T �����X����:1 Wc`f<P��DjX=K��4;�N�8D����ڶT0��C�ٗ	�zߪ��c�v�����&��M��>�n	,�8�-���EO�<� v�ng���^ڳڙ ����l���k��v��.0��ޫ�����#s���ϡ�	�Jd3ȥ͵)��
g$ۏ�[aI��[�m�|7:�	�h� �	��FpNz��Fv�WI�mK�*s��[uLd�ͫ�B��0q4a��c?u1M��vv�D�$U�P�dG; Ց�i�+�B��ƶ㎴�/uV�����UJ>\iѭ��C���͖;l�{�KQ9���}x&ƭu����E��z��G�p�&�q��K�5�ǰLt���Au�s%�N%��xW.�>d�q ɲ��Ϳ���=�Ğ��*c��!qN@>��T�Mi'���=<����!
YfO���5��3Ǯ<u�(��ȉ����#��	�96�Ӊ��4�g�K2�OX��Z̆Z�I���8��˛��t����򬦤	��P�&�,��ǶJ*�'\�k�g�jن>�|񦓝���e��O�{�`�^�����l>�2��N.��~֩4H1 ;����)@����-!(��?.�� >R�'�Öj��걶��bLr�w�V��Z���w�>������뭹�9|��t&P����ˈzp��o�M-^e*����~:I�"�֊������0[�}7P�6g1�#F�w�YK�ݼj�y��ا�/8�ra��(���~�܇��"��$K����P;�'1L@��C�"8��)�� ~�!��س������_��8��a�3���bQv!�E붼 �tD�o�#�+=H�l6"���_���dH��C�R<�z�[���u��/�B�U���6�sg0�.�Yh���_@��A��:9@8�o�����te`-�����͔�&���B�!�	1o���"|i��|];�qY�ՏK+�}cL4�@WV�z�0XM��7ȱ��O��f����yr=�ٸQx�� �P{[��:{��E�6<����l�~��ė���_���6�	lk�D ���D47�E��5h���֯�bƢ�zәovO�-�  v��v�_�`-��r��";?FЋE�Ky$JƜx���0�N�Z�x�<���L�O��dpi��}��1b�����Ϥ���-3n��͔9��*�������#��#����j�uA=�)�A𺆄SN�Vo�Z`���p��ΐk�9LAy��u�O�E��y��-��B�.��}b�K�Z4_�x�u�V=�����I���~�9^d�#Oo��މ)W�L�pe��)�W^rY"�0^�߬.�?
`�@�,����T�nR�N5������<(�������[��m(:"՚�pal�fH��$�F������AC�_�������QĮ��b������vl�t��G4��q�`�t��Ko�������f�&�2��<v|�7�\r��s�!~+��W��
���h���0zY� ��qh������Z���2�ࣦ�l����^��7
�[�p����M�o*���s彴��Tv��ZEmc�5j�Ig�9k�W�hw�/�%�0Nr�:�r�Z�;
�o9X��YK���.�ѩt��Vؠi՘��#T��2��zLdm<y3Yj�V
X��p"�6{��w<�l������>��������Wbp_U��˗��x�b[����tnp�<i�}.�0���\Ŏ���H�֟Y!R:ꂶuW���9LՌ���D_�T��U���j	ܛA)c��_uNd�I:�T�ٟE7�@n�!�m����&���c�tw�P�v��n�Id6�hӒ&�<�ϔ���D؅���}S�
E�y���e�X~r��`@p-9]�j��M?���3�8>|�e��E��2�g��H0T�-&M.�,0$�tz��(J��˻^]��/�N�z�w󞔗��MKo�d	ễ��2��,�LdU��*Z��B�(~C����\�
(��\�?�>{��9�"&}�1C����ai7y&h���B���-Ep͉ߕ�!?�4����E�}�SYۀ��I_�3>����+�o�XEJ*r4�R����i���jZ��в�������8���a}���*�֦7>#�����!�0�@Ǿ��4��a�
U�DCM"#RPL�-��+��7��,^V��{�_�T����.MrA[��S�(I���	�ʣb��{\�;<����׽��	;���>��
sR�oZa���hf��(�"�����b���s�IX�)�U��v߰������M���V*&�m��u�n�dűv�y�Ą3���@�����O�s ���-��M��>̩���e"������ji!�+I�([��{��"�`j١����j������aV�W�JiY�\��Ⱥ�DD�@�C�Ë���j�ê �V���'s)�_0Ca�]+�f�r���4��p��i�+����8ۉ¦D}ﾈ����s �%��=��fb����]�(�����
����Me�������2�y��$�t����m���n��Woz(����&��z	$?{���O���3����5��z�����ȄR�$j�t�>�{c�O*��\��J9Em�$�z&g�N%�ݔ����9�ckL*��f�笥
t�������LO�u�ܦ�����ۉb�J<��7@l��hIZ��<��R_&��݅��&��B��=���Mr�ev�nrJ�Sl� g�܂�"���ܿ�m�e~��8�t�o3��X0�Zp�N+D0gI�\�_�5�Ar�/��WYh�L�ǐ�a��k���T�ց��?�}?L��=�vj$X7bS�(��ݎ&�"I	%0�y<�b�6#Į����7x��]�f��w�'A曖A�w��jbH�CVCaVS|ŷ�BS������N�53*G��p�%��Ȣ@4̱��-:D�$�&q>'�z��Pj!�O�W p���,�o"$>�yT��̌�����:�$�A�"H��ekb�M�1�_�槈�Ogw�r)�{�Y"���ǻ�r�X���g 惟�*�psGg���b���  ���z���n��T��t�!�3�c
4��:X�nz�_����9��S�e���d��(ܫ�t���;vټO�K���2EmD r�';P��V�(p��2�W h#;=QR�U+���WZ׺�@������X�z��������ꅯF�$Q�P,��_�ĝ�\�F�mU	���O��1�Ż�5����4�_���NU(�>����6�Y��QB�r����_�ս��h����I��`���C������D������Ǌk;�]/B� V"�Wd�WmP�S�V(���*�13�.�V~fP\���=e�l��B$@_�뭊K�x6ˌ��Wӣ=��8yPX�4��;�)����M�uOޯ���6�,�)���ֲM����H����[*"vh��6��'qn���Ġ5�Z� �&�+H٥K� ��^��؏�K&G�����!�$��$]cv�eW|7d��@|�#��l~�ZG,���];o[�4�����ni���Q���co0����y�X�XY�da�{�'hmAG��H�fU��x�\eV?u`����oR���[s��L�S�C2<鎱����Y���Q1�����Ux@�.�%؁!^Ǻ&�Q�m��4<ο�:ۊ����h��K{FA&���,PN��}ͫz��9Gػ�L���-�(L-�s�2��*=���=V�d�����]���3�46�"�z��v=v>@㫤#�.MM��y�Mo&砝��u,��d�1hp��miz.GR2C�]#�4�Ú�3��2%�#WlDc>j���U�ڰ͐�<o������7ypA�
�W�����g`�}�c)���O5���C���i[�MҕDW��&�y� ����u�	���� �����[����m;x|h*�	��t���� ���y�WPi^����4C|�x���i��yw�[�]=b���(��)rW��IN���ٲ���-
����iJw�r�"��V���y�RP�N�H�ջD���9>�&@��8}9�Jҙȑmzg>)bpu9u0yk!�,�Pk���3B�?v��I����W�.t���e�3vX�z��K3������Ϙb�3�&���d�C����rOO�.�7��`=&����Bй]݊��i�ɫD-��btV���2�ᯡ2�^��g��N�8	�#�W�	��'#�Kf�!q[��>Q���������}�	m���$�j�{Ɂc9 }BK?�X�^YT�3ט"��.�+j�%�`��%5V�òG�.ud�$����ȸKWp߾�<D�����G��S�� ^?�����S���o��� ���@.F(�b%�p3)2�i����Czx�f��ȳ�=|��u��]0���B��X�L7��Ff�b�H^2�G��T��γH�|�di1��y�k���
K�G�̓��q~6F׮��MGJ��l��h�,�0ȣUh�}]�.(Rk�e���awDM�1�D��'��G�[�\rGTf��h:5�M�M���Y��{^z��hU���5�= ��m%��΀�)�4�5�,�JL�;:���`�a�
ƣ��?�0x�>b�Й#N ��Y&�����8V�QU娯�6�+&��o�bE��7{��Ee�e�SJG>Jm�_������ˌ8Ru>���Y���\E���Pvrs���Y��^wy�>��jS_O�â���HPjkHD���Ƭ����U����C���P�h�o�����A�����A�l稽J8���}�p)�$����#)�[s�6�4�  ��v��2�����4��=?L������.�H�>�����|f��g�J�sk����)CdQ�ԉ�C!�4m���g�F�PM���h0(T�!9�W�lf��*� �ܯw��?��^��1�'<evބ,�+Xk�I{X��	�{�N̔����]$|�ZX��5Yi��}�;��]���#�o��wm*�q����[Ϛ�fG����{����4��c����S��CSݞ�m(Q���B-LJ�7��=RK�5��&���^��e��kq(I�y�m�ִ��`9���8��jd�8��}��������^�x&4��%�H odT�2��:'��K��@��������>!]��A#6���l�}�:�rb���[�`$�m��
���n��� �b�����G�P �0:I�~���7��h.4�s��5�1�x߾?���`����A�@�<W��w0L,!���q����9Fp�,eF��] �C0%I�O�\x���J�3D߅EP:�:h5U���Y1��%��l���W�
~��/fa!�O���Icv�5�+��?rvp�I3*��aT.B&�0�7C�A�%g\�B�Ë��m�o��/X�[#&��,���%�{[h-�:�{/~�Hz��߇�4܃"���4&o��p�>U(�86/��!s�#e}�I�1P��e6?eIz�틹��N͵|y�טt��Ql�;�~'�� �a���h����N]/�)J�ٿ[00������PH�řYqqr~�p+��5�C�b�0I�����H��Vb(�\�S��z�1��<���	���<��Pm�z=u7���B�R��G�G��_�8��qnߣ��(|aox-}�&73�łE4�v_�o���x]������ޜs?<-DCS��x�}�����@���͊�[��,��~R�֫�b��R��Cڌ��b�� ��V���I1�� �t�8�������؍���}�`��h�Z��ej�y�4�&-@�=��1"��I��@8H����)�}��e�%��I�@T�j�DB	�1n�Xo�K"�+/O1~�(��ĉʽZ�st?��(�njS������åӃ�����V�"Б&�0K�S�\�;�U��G4����U�*8���d���b���R
M��p�}�S���i��Hw���G�
�ԁ�̶gRm�6B
` tT�Ʃ*<����@���g�fy�l�1�^�,�OF~��0sk`��ܛ��Ʊ�'h�����/��q�i���x�o, �_˺���Nti�(��i^�h#'!z�K�0�e����U̻�c=�ՙh[*����<$�!�V8^3-m_���1�\ڮ�3��g���W�F�M�Ny��zAtG�.� �����pߟ��(�?e7���2"R�d�|�72~:����<m�nH��־:����@����/!j��+��ml������s���%�o ����G�3+t��%�m���Md"��v�^Wx��M3�K�"�0e/���ʘ]h���]sK��o}5tj�8���8�bp5�$
�ň����a�GJƈ����G����J�-Xb���U
�	:��&�K��2�p�V�y,�Hw�>P��R��}��9�����8^�*��߱,� �p0�RF���>�r8Yp���4�89�UFV��YB�K�G��&"���'�[��w�m���I+S^Ӄ0>K�uz-7˦%��蛴f �yB���.�Y�H�d@@߯�r�������M�ђPXɹ���O��ҭ��S��g��I�J��8�$E'�NԞhxI���x� &-�H���%�s�p�����خ���)�w�V��"����y��������n�3�F6)g-�ě=e ����|	���Z���>��x�<�����X�!@W�
?�̽hHH}/&�@@���в�'��[}�hWi
,o1�yt��$�O~ޔ��G(�rg:�6�oO_�L��s�4�1�V�v��T�"�(�K�+PLY���"!D���Z�E/�S��]��l1*nԲR�ۦ�D[�fJ��Ք*�#�Ģ1�� �D�{���$
4��~������Ų+B��^	G/F����f7�Z�{�*�~���%�]'S�Њ���]��S*7���J�#��� =��*�����ںT��$���Wdxn�N�y��~�X���~z)}  ST#�v #=1�mX_:]L,�l�_1��>�8��đ#$D��Rk�{vt�])��h�����o�ك����4������W�~U��G���m)�o6�P��2="����Š�d ��=��_kȕ֥�x�Io'�����F��*�Bc��sY���&�p=_@��r4l5N�U{�z�*7���_�Y-_뮝�t���� ���\Hr#S_%`W*6O�Cv�T򭱋��ČW�3�vRĔ�wZ��k*)iپС-Tz�i�{��DB�N�JV(�0p��8X���R�_�ԃ۞��ۿ�
��ZW"/���ʙ6qo�N0��އ�M����_d��㨈C9��B�x6�M^ F��d��LZ�>�r4�v C���>��n�hNȌ�9oEsd��f����B�oQ����;��~��rpab�uH��o�G"�#Gx^2�gdvC��i�s1��H�B#�v�>��:�dt)^{cYP2��0��)��q�c�5���?��x�eɱ;~C���#�}�0��P��EL��ᕘpB���1��PҩJ���BY[z�u�=������3��7� h����f> k}ѻQ�F��+`����Y��Ts#('E8�SG_������)\)��u���s]S63�E��[ژ��]s�.�Ȣ�O�q򱕔�	[^����� )�P��8��
����V8�[*�nk��X�u,�nDE(�2�0�&\�{MS#��>b>Ǒ|��*8�l�s�׃a��i��Ow��~��C92�scC�����e@%�W�g�#Ky�d\R��`6���6�2�.��~���c���&����;u��p��ԉ���}U��� n��-׷�/����c弍���譥���ZL�ܱ��C�]�B�� �"̼�|�ܿ�?1=�% �T��D�k^�q�����(��=�n\�L�w�u ����D˔��O"6bܸ�@��3c��'4�K,d�����&�]`����8w�C������&JE~�5��4k&R�Z%	Iˆw�5�c<A/j��	����b��H�%� �%GTi3�k�x��su��ؚ��qJ0X�����]�	���-��6�,1w�)���D>\� ����[��J5�V�sE��2��/��V�A�o<O��tH�@����CCIE�:�3W���AY
�Ń��gINK���Y6���_���L�N��5����\�ߟ�ÛRp5>�p՞���9�C8���n+�D�%��E��
e�֟�Gs�Kb���Ho�h��EY{����Hj������h*5w�B�1x_�ǽ}Aߚ���i��$A��1���E��yR%k�>��G+����q����H��{�+�ߝ&�*��=je�gCm�E���۲����Vq�0R������:N����U13�Xx{�n��p˾�6��rN>4i�5g3�9��D?����тp";�jL"p@l$K%l���b����i��:���{�<M�����LIz���+f��dV�#���:�l:}��V�R��Z��g'r����-w�ǻ8�б?�:���
&���#"塻Co�:����"��eq�֐��-^k}�'
T�� `>=X�w�B�s�.��t�6�^�f!�s�T�D�j��2�|�P�[�[�+\��2�=�	59ڞ|�T�Ň#]a���!Q����.���a�`s3A���Yfr�}+fR�F8����'G� ުˎ��^�y[p���~~���Um�}�Y˅W�N%��a�k��&t�9Z%��V�F����'eLC�!`|3��5"�� �rt�V��7��a��ִ�.�e_�3���%l��q4���X��3M3��;Ѭ8ҙ�ĕ��[����&�,�+�؁.Z�_n��A�y�;�g� �� *?S���t�d�\(h���e �ƃZQ�6��W3":6�C�?��0��4I��P��� 0B�_�).��@�-�H�XC����fA/k mŇ�1a���i&��;q�%V�a���8�Ar�����p�v����;�?M|�\��9j!�I��n�������DH�g:H|���*,��V���O.����N�A4���H�����z5z���y�oH͠��!�ik>���!����vn�7������qt��U<���/R�h5q;�@��}-"�����em���t�|5�6�@g~�:w�~�cj<�l�`�|Q,�:��Hb�F��FkG��$�Z��o�H%P�4߶{�A�0#(<��(ߧ
�޹���Ʊ��D0���#�o�,nK*�<h�..c��s�W&=6�+9��v$���L��4�I�Z/}S��x��M�v'��%�w�^�C�iY��m�*0&���d�9�rDؕ>UL�����bŧ\l����+���:(�����^��h/��GL�Ͷ�����ս�����G���_Ǵ����-[�j�!� ��+��*E�S����@��I�����F �|d
N��t�o��:ؕ�����7�(q�>ǖ ��z!�֟�����fў�r��W]��.��\k�+��Q@���O�R3	���^�/�
�P���] �ކ1�}'Ⲏh�>xri����� �""��%�t�
��zЙ��..��k��ٵy3tclZ�G}�)�p>����xRޏe���t�6���PR�zYs3z����v*����	�2=�w�4���D�)h9H�q��Ry�������ÙR�`X+���׭��l}���������q�>�#��R��?�q�dwk�1�h;�p�t�g�"��OU��axd�t�� V��$&�D��	��vP��F�1�S*M��� �њF�~�x�ٓ��ݰ����I��Li�q\�X����-�z�P���MJ����Yvs����h��h.~�Β̑��ͼ0I}�t>4�>��t�e����^�����''�u��$I��;�sK�-dv�ej	I�V�,��R�!|V�4�e�ׁނY<��[��vF(���z>�5vG�,4yE�T_(���8���ފ1D��*?{�ӧ��#�}܂21	H��z�~�]����ik@:�A�ܜqI�;kyDS%�G��8��� Z�%�j�g����;X���??��ڲ���)2%CX�r�͔=�oH�
^���&z+�[��&ay��h�/���Ǌ@�b�4�񕩩ӹ��lf�9S���w�p?3`��P3l5�ǟ�K9P���(��x�F������
H�>=�9��J����@W%��F�Ny��OQcNi������`%�B�!�����V�J�X�C͹���#��Ϛ
�5*(����`P���~l��]:�U=NY��|z�L��1���[#�0��0;W��fo�6���Q$%�4���6�o��$O��:�����H��b;�<�	��~�d�m���,��q��6�	4g�K�
�_��;e
]Bɔ7�ʄ�kӓ��J_L�~�Q���BF<x�h��졓�.Zc�����h0��;q��
�kK��(�t�t,��;c��h��	v~:Y�9��"bt!����A�:^�y�_�:T	H�����d.M����gE��|y�F�/U �%T��r�q��e|�6�Xic3���,�GR����@,��R-��\�7vI��\P���rC����u�� c������{ �uw���v򠹩זּ�!N|�H�4�\LC�
}������io�Q����lo�~��<����<B�qV��4<9S�F@�����?*�����}Q�\�ũ�z�,bGu���&	he4P+�d�\��͙jQ���O��ɓ-���H��(��c6�x�6AX�/��g
���A�7��򻼬�1��U��LܤX���n�s�{>����� �ճ-���j@@(�"\~ݓ9�~���Wlt\�p*��ECʹZ�Lm��E{�x$�l�Qe�U�P-u,^��d��i�,,6�g�q��F�4�pE���]������m��`>�N�i�93��gA:j�i�{io��u�5����!�[���ջs��y�H���3���%���N07�v"* �i�˲(��K�pqw.��d�,Ґ�_O羣��0eA��g˃�_��&bVj�GU}B|�R�T<��X���q�V������)�ز�i[����ќ��A�rF}�&��gqTҬ�ظ�>_h,��,��5��ֆ�-��y�^�0�os�H���T�A�C���:�͆�(mj�6'[K�c#@v��^A����j�/&~�r�@������<��+�����F'�8�5���u���Cy� X�?�7�� �u����{J$���*ԥ�P� �.a86�2nVL�Ʋ��I�<P�LxkT̤-KUω��*^W��l��ofǐq�3pD3�W1�`�Y|�H�'�3S�(�����F���G��ƭ��/��l)R/�G �+�TDb���]�|�
�E�ȋ~��q&�D���תr.�*����WĸnM�7��Y\�s(��NO���F��/�mފ5 �4�}umR�Fw^=4 0���u�D(]℆����������e�B�r���E+(�Ȟ��nSO��*��A�Z�W��O]�S7��~ 2�t�L�4|���>R�:b(�֢�-?�آX�3����4�O��d5��3�8��pW�����.% 4|����v�8׭��F���=�z�2Mo�o&#wܷO0�+=��n�0[E&�[	�P����t#���Gh!d��1j6Wr��2���cq-��Q�Z�l+/O�F��s�Q�Ĳ�,�g�I�q�dm^D����|��9ݮC��&�o�y�~y��BR,ƻ�Jk�Az#��A�Љ���C.w2]�
�\�&��{�W�+IL�� �]2L����)FM�Q`���1��u�RM
��Š�
��f����Օ<EE,����wzR?Y&�^�d�ݯx��o_�s��x֐�P��O�qIc�&��r�j�iþ0*��EW��6]D�2�&^Qy��2ԋ[}���-Uڠ��6y&�˕��MF�wv[��)���g����'j�X�q�S~	ꔵTt���>9���O)/����@j�^����`�Cx9��\C^ޡN%Y�p2X�"�4|�]xb��+��צ�댿��D懦�ߨ�����z��Fn�l/]�x2�q����_{7����8%�&nq��<.&������S8�> ��y>��S�9��qrD�� �U\����\\$!:�Ħm����"��CG��@9:�� ��4��ʡ���[uh�y=J�4�VU� Mp໏��
��������ۋ�h�W�i��!�
�?��«ʆ���n�c�������$j2�����~2��E���� 40!c|�]��I�uD(]��c�2}Lͽ�R/��we��ܚ�񸎋
�}�{#�[� �Ǉ9NMgTI6�<����ʇ�&�9*+RA�+K�''02�[i�3�ܚ�?*���b�����{aT���l��蘽9g�G�A����pM�f�K5N�}�Tǖ�
�b�'{N-�<I��'/�XG>��ɗ�=ԴG66M �����oidMW��,�+����YI���^������t���a��<��k�� ��۲���-V|�Ĕ&p�vw�c%���Cv�:8���zp6��W��)���ְP���M�}�k�.3�_,�۠�M��+AG��+�c
�y]� w4|�R	�q�ߍ�+�e���ݵ��L������-�JhVN�,J$Ľ"y���`]R@82������=R�kQH�+� �W�<q�v�]�i�S�2��0��b?���An�f�]��?��'9�F% ��{�G�կO(WzS_�8��n`Cp�6I�i�W��b�����;��I�=��˭��Xת�e�q\�(�]����v�/V�Ӷb��Np��k�Gm���CR�aw]|�����44,5�F�o�����1\E��Y��md	g{��ҡb�-���`[pf:��YaD}c!�C*���{�p�b���Ψ�e_��������ð��xM�K!�ސ�,�(��yJ����i@�zPH%j�g�/�a\��o	�a;���҇l�?(������P��_yll-T���O�R�}{'֡���iaQ%_����-�	�M��k���t�/���������t�Y3���d�j���gwn�_��¢ҟ�vN%y2��pK\}�&HeI��-���bfU�Y�0)�s]�`�� 9�#>2⁲L��I�~*i�rٕ�����@���ל��JWpt� �|A�<qk�&/hm�(�������d�2f���7s"� `Oع��}aᢜp�!n�W4N�����,�W�N���' R�8��ܷEbc�����6xga����e���_3B;ƫ=tH:lp_µ���.8!����i��l@\���'A�Q?�.��U�=27I���4���@?� ���Q2�	��Y-�fNڻr[Ca� )�j���F�,QB��8�Oa~��@��$)��OSze��O�#����i��'�4�Kh��e���7F%2X��ݷؕ:˞;�7g�D�}�ym��y�W_$��OR���%�*������њ7����M����Tc���o>�+f�E'RS���iQ����y�F�0��t�Ԅ׼�d��'�g���*hC��
!��`UXжQ�;y������*!dZ�@or��}:���e�D���*+�ɳ�`}� ,\Ï�l�l����8�� $K����w����/�����.RD0D)4�Yh@aǸ�����0�\�rc��x�j�����de;K�q�����mm%��r�I�7�����N����ٝ��W8a��������.����z?!1��$*�О	8aV���˃o.�E�"�g��𦪊�����Z��,%ryk��>>�e�!O����)��辳q�8��2�F;�k#Zq�����:����_@���+�#�<��8��*>ƍT\���YT�S~d��������ڼ N�[c�D>ở�f����T ��U��>2��=�����!���
�r���/�.��^Mގ�����������݉oo-Qխ(0�j�%�(j:� ����B��Y�9�h�d��	�X�3Ō�w�	8���۩ױ���`�?��40 ځ�`$ӈxܦ�~��?�BHd�%��y��^Ȉ��6�ңw�`DeeXU$=��P*;�vCƆ�D������G?�*b�
^!&�$s_��a��0�N�%�2e���`y�	� �e|a��H�%�B]F,x�����@���q���svԟ��� V^���݋��U
�����>K�ac�@�s�ʨ)�s�D��˶�� ����p[hT�q�6�z���5uǜ֩��B�9�Nx�t]VJ9F�6�`q��'�=�UF���kes���Eϳ����ͻ�{�p�Y���nLz���山='D �@�塖g�i�u9Eu�Y�G�D�m�����#�M�dKѐY�v@̥��C���e؝O�R�"<f.^S���~.|�����i�g��pF �͒Y�;����3�A��+�0�ns�>�S���]
y��������������I�B�U_������-蕏!]R8�FM�D��B=��'�^�Up��oR���{�ȴ�v�-I�k؀y�W������
���L�9���e��,/��}�0a 2E�Ɵf�Q@26�!����/ 6�)E�`�q  >+F�̵��, Es+�M6��Y���vhƗ��^t��=u���Ѓ�*EW����+��D�������ܬ�v91��������a�?|��~���*���)�e�A�''�g��H
�1�ՙ��ۼ̨a;]��@=�x�e���J�V�\�d5�Q��9��-H$�8�G�Q�uA&���p޵n6���o�G3���NU��~�FVfr���[?�Wf�+��n�y����J�P+���������Q���d@�����q#]��ڇ�ϻ���%T��$���1v$����t�`�9��+���[�6�!9���o'�}xkS;q.e+w�G�@�_��Y+������(U���υ���Yjr���(/�I�{(���ᓃMl�H>0Hz>���uK�����h��aI4��6�K����6L�E��U�5�Q/���wh������&�(��(���_���ڂ/C�	=8��@�`k�q��/.�	MNڂ�8��J�** �{����ي�
�Z�b��7Fx�<��(�K!�9�1�P;�Z'�L��"�t�Moϋ�����%�=��k]��:��4���'���C޻pO� yyHT����4���Z��Q�*b���*==��eظӺ[}H�0���\��N��a��i���we�B 2u�����d�GOD�M{c{���M�t>1��T��YX�ʰ����//0��~s9�o!�iν�,c/��>����^� �J�;3ϣ=�����qڧv�%
�l�j������ǯ�9����D�����G�E���"� ˺��e�!i��g��lit�����8���I F.;;��.G�O����h������H������KKQ]t���n��ӖT�6�`��V����^u�=����O�Vi8�w#�hM���K�6"�ռ> �6)"��Q,�{�k�Ԍ���Pd{?i|�����J���=�S=�-��x)V��M�ai:�s��`pƱS�j�V�pĲS����w��k]u!'[�g�?��WI��	�Msz��N��4����Y�y�vή�#P�y�Œ����Z�T^�6�6:v��̼O��K���a\�l��#80��)�5-��:�-�\���Y	�����Shֽ �.�8=��e��	�r��=�OQ��.���Ϳ =��&E��i�����f��:�/P�}�g�i�m��Y2�0���.(&��&M�|RR���Nf!k�!_���o✾	)׌�r�A�a�6� ��AX�?�&�ы�� #a�}JJ#)��=�h��W�M�ٮ3b2r���[
z�۶I:M����ʓ����Z�w���yݜ��Gh�#�h��m�n���|k��5�8�SJ㱣�ȿ�ͧ��(Z��&����E�z����l�=-��7���Q�Gⷈ�j�r��_a]�P������%�[�{�X�U�e'���?9
'�6a6���u3�Xo����ۋ�JMx:���d\�@�򿕌l]�M3U�9�r��<y�Y�y�Nn��Je��s�}2��R����Q�f��|c��߱8L_ʇ��� ����;�u�sa��<@6�L1� �B�t��Q��E��x�ef�'��f��,�A�a�M��#���"7پ�I�bi�8�������¸��KҚ����K�/y��᧓��}��-�i ��Nw�d?�����5�e�7E��c�
{��&���b״Z�n��-�X��6pU<�ĸE�j�NUL����Pɞ訩t��U~=D��5���
�e��u��򅜱�/�����F\�T�1�zύ߶[E	���u�<-2�C��e�v�N��L�à�ِU��G?=���/'��!n5��5��F�{>:���M�|b?laRİc�V��k���;�J=�v��zy�C|oX?[��h��Y�K^��y_�<"S@�%pu	|�p
^ɭ������v:=������:^�|�/~�/$E�����9@{D���.Ȣmݥ@*/'�^ߗ�ZR���0�R#�������(7�9�L��'.����3��Zͅ��F�[(~E�����nVn�=�<Uћ�w��.��C[��O�=:$����ꑴR���Bb>l���}7_�gM�칒c�.����we�	}��O�>�G�\=��.V�C����ʆw��:�FI)Έ�K�r-%�'),�8 ������l�\yk����	�zj����:�i������	fO־���q�	�,�3"tW���8ԨRO�8�F�}�e����y����'{�h�o�,�8�r��^����]��������=s�̩l�YK�حg��Tˮ�7�ŋ�{}���p��[�W�[N^O����޺�G*����i�[[��00E�x������w�P~'L3Z;A��!$O�G و����r�O��d�V ^FQh^-�'�c�#�m����.���朌AOXoҚ�h3�@�<	�MD�O8�[�k^�|g1,#Q�*�Vo�B����K�-'	 S��m��b����ºF�NJ~%��.Щ�1D�v�c��J�Z�Sȫi���b�;E��g�Pۢ�zB[�x�Ůu��Y�����qLc	鼠�4����}�ϋUCx�EP��i����/�o�^d�s�0�fܤ�<��I�uEאFh|���T�\U������s�}K��;Od��?��8f��tZ���,۪��%���E�@�yE�gz�s9p���կ�T�,�0�Un9C�I&ł�e�n����~�Y��^�$���&�^9쑣[4�>-��gbU
��8q�&�F����:�Y�2��Q�Ƽ��%Q�cm-��D ��ӓ��� Q����\ug��sؗ�9C��ԯ�h���U����А����5U�����x��d��L�ak������P��;&�CO�li�羃%?�R� k��Y�������Iş�@<;�¾ԩ$Z� ����ZP��c��֑��#(P-nڜ����(	���2��52�xu���ꨲ��ev��R�q�RsZ�"
�E��o�a.����~�Vt행Di��[T���Ύ8nQ��䢑���"]���d��G��RΖyxD�������i�=��}Di��`d���ͱ��~|/����6��r| H<���{E���E9��w'p�c�n��8�����}=C�0�#M�@еb��$�*�;�I>�M�E��)~���st�#�������,F�F�RA��7�~s�@-c��Mf�v�u�v$�E�ww�>����IlR�d�(�8'�N�bN2�@$����|Z�*[;Y[lu��s���tA��פ�a��&�hZ��Y ^]޾����v���6A��.)�f�W��g���uT��W�QE���q�=����^˒c� ���d�9�<�ր+��|�!��(H����4�N�q�=sE�y!^FS2	2��$2�!�H����dcFYA�����L�y��T��.��w4O�2,X�+��?�a�-�i�ޭ�"����1묉YXAw�r�30CNn�̕��ڣ@��~ �-���Oi��,�b��C����6�C跂���z�����U�OY��R��^��Shj`��i��u�P���@cQ���/}i��q'qc����A�L��΃������WԧT��t���t��ۥ�P�;��1����-K
��6CȞ��AkZ��������ݠ�ë���f��^͛Z���������:B̝�#g�1ğ:'3@�o��* �H�;�//��O�s��������z�&��6xb�;6¥:)���#L����P����k�����
�yw��2�)�ay�ەD�D�%ڼ�'��0	&�
����n}����rpՇ8Z��#��
 �Ҕ�ng��WW6C4Է.|4z,a��C���]KZ��Φm],Y��[���O@f����	�
��H�{2e$�,�L��_��)�*�H'�=������]��q5�{PL�M�' T��lt����X<|�
E�1�*�P�(��ϩ���3K���>`�|�g;��Y��,ۉSC�o����9{��zAi"����9�
�&o��:�oÕ�sI�S�5s���5��v�b�~3e�p5~��&bqt��#����mv�p�'��G���S��L����F�g��������i��:ܧ�����J8���i����$���+��h�:0�t��>.R�7kSld�Y�a��V���Z"A)�GZ�ژҵ��̀CD����f`	���Q�_����u)=�[W.f�T��w�3���o��ͪ���x�)/Y3zƮ����b𸯬	P!�X�뒽�!�6VC�/�'����U8�P�Or|�/w$?�̾i�^(�"]�ѴTD��К�����wlB��[�}��Ba�@}������3ܾ��\bq����Bh{rܟ-��X��<�@��?X��R���r�^H�8���O��&T� ��%��%>���u�B�6bmش�������=:�6��/Ó��+y'm���GI�������]�~nUb/�{��FQ�D�d�7r^ �l��w��gE�bwt#�,�wx�_�����!/�%�u��'�D��D�R�u�\ST�m�	��A}�E7���� h�G��]"뛬�|its�>��!��C J3$�c�:Q�1.[#�#�҇�<��դJN���n�9o7�����T5�˥��L�/s��>�rԔ�t���q?��S��1������gL�K���|�Ş<�='C�J
�:xTD�G13�(���0�Ab]p�)�<� 	��%����>���ը�s�{��?��&r�8mԥ �)%c��_��������M2�jY��.���EH�~Z�H�n29lUy2~v}e{/����W6��\��@���+~�=�&������d�o�b���0���A�n��@Q��QK?
n��x�n���*�.�1�!��棇����RJ�۩<�HW��*�e	K縷�����(���я�0�-�?jDLO]~�d~"2X]��aA��p�mC�U:�����!K������^��θ��q�-F�50�r	K�U�a,�R|ʎh�����T<�k���/�觪 	��/|\��\���gC��@�,&��?mn��y�ݵ#N��a���2�g�J��C��H뺇��L�	���g�75vC�U�L���O<�(�! ��Ue��Wg�DȎt����G�U���������;��̮�9$����W�H&g���ؓPy�rHZ�.c8�l�/�b��}(͚���|%�'�V�3�I<�)Y\�c�HHpvQCF�C5�p�>,�]�ć��e嗙N��o)nVPO�}�9N~��B��g�xк:��g
�~\�:1�b��J=�<�%�AE���7�j٢
�lP�X���/:����Q�D[��jԲ��{�5d�[���7qc�r�I�G-�~_��e:(HG�04ۚ�,�h�n�5�/�U��,dV����i�H�:7Pa���b�����RgUYmSg���3��)o���lf�?����ݞм�t��\z=`Eh��69ޑ(nho�1Nuo���J�6c�fܼ��<�iV���)�ă<�9�-�|$Aw�C�d����n� l�|�񧟛�xĘ�Р~Ql��K|J~z�f�T	C/y�	��P̚�sAR��),����Ϙ�a��Ы�P��蟾���E;)K�ȏeB���۵$*}�>�|��Ҳ�VPL6Rq̵��s��ͨ�i�Au�X�rXܟ88�"Ʉ&=�2=#4<�$Fe�1}h��ӌ I�.5S�L�U]4}�fq��E�Be+:%���2��T���[ֺ�k�?~9�o�ˮ�>�.�xv��*�Ǖ��2�홯��|BZ���Ey��d6�������8�YR�q<}����.�v�}(J��7����W׈�4ze�F��^e�p-�un���~q���-�XiÉn�S��p�I����=5i��|mhg��y������Fe�"��!���1E�6�%[�Yf)yo(�{0�椸,�7aP�P���f��B3��YnR��n�A9mױ��U�������E=m�i�ɀIp���O�gL�,���;��3+�Ё�
�`�bUF��].�rk�̸ �G(��s��ɽXM�	зtmzKn�� ���a�Д7�/���:�oxQl�BO�HX��!s�j���-ăP�������Yױ�	fʔꯓ�gK����"00",0ҿ�Ш{��`?���QW��IkT��#@�F/�U��w����N��%����=�(M?�9}Zޤspǀ��YLӅc8�1"�9������	�<�J���m,QH�vYf\ߣ�S">h|�|�̎�i���tݔap���I�qHR�V��� $�șsD��ļCK@ ��ό�m���r�J�<���Ee��P�p��x�	ݪ"�̅��K�[�6Wc��P�-E�7�ד�֏p�5�������
$�_��ϔP�B�BPsd�M4�^:�<Q�G�c���Z����4�ƺ�ϧ�?\�ztq���z]R�f⒎�m�p��3�7�̸�`��D��ʔU�u��3��a���L��=f�W����w&"�J�rc0��|�W����H� :tl�*`�&��jbE�y���GFm��u��Z^�#� |łt�߮���f[s��Zp�61�V�΃�4�'�$�W��� g{f�?��f�l�DUn0���yds=��m��L�K�d�*jR�ԙ����@�Oά}�)K 7O�������bhJ�z}��|�iƸ̩�4�E�Xl�e��T���|_��{3��'.���t�Ia�3�>�*�3��M�Y�Zu�{ݬ��;��
N�4%����cSF.uvC�*_�&�m	vc�&V����ի���P-z�1�`q�����Q���)���of��|*=
v�Էu�b\���g�C�y�t
��D?XtO����Q<U�$ށ�~&�y<zwaۺ@�%~����TO�qx��)��n�t���
�CN�s�A��XƿsΩ Q�9��bnr�E��L"���R ��L	��Uߩ�?����s$�;?m��XK�CN����^Y'��V��4!�q�V���땿�8����AU����>�kpjWT�"�}�g��"�w�G����B�e�p9�� ���S���\��Gp�l�p����B��j�U� 1{�XӅ�S�Ml��M�Y�r��DW^�������K���Dv�M�� f1E��v�@-w�/�&(�ہ���`ɒ�����I�rJ)!TET�F� !`չG��P��R#e��Γo]��Do�G�.I����qne<�yw��AX�٫%l^���%��T��4�,u�j�\��9�a�JkP��>��;z��W�T�$h��O{�7߹ ���_搴�#�>EN�!Gp�ԩ��|mx��xG���՞�ܩ�[�o���t
��_pe�3�[/P�!�MN�����X�f���n�,�hԽ<N�Q\3y��疄eS<ó��?���e���!���AG*�1z��_f��R�J|�M�Q����z �M�?�c�̞������Ĺ��&Fj^.�qJ:����TϞJr�)�����~�ߔ������!kw�p+X��)gC�I�����Rhq�iW?�ܱ8��\:�UV�d�9ѓSUJ��+7�m���}@ ��B��a�ץ-\Ǵ��sDWH����&|Tl�2C��;%���`�(mW�r�goо+V���Q��hK
!��N#:�і#�Pb�m&��:�,�=W/����i\+�������a?^�������Y��y�����v*�Y����'�P�Ͽ���b�b�G|�ß���S��:��cR�,�t�?OXĂH-�V�C�1h�'t`-�.W'���3&I;��n&�/b8խ�E{�w�]��Ӽ�[e?{�t��@��8ک|�a�hR��Ç{����C*��_!��,D�U����4�[����3�q�[*�1ш�v;�d�v��r`I�	��ȟ}�w�a��vI#|~�u$�2����v�--_]ݍ!Բ���ToA�z\��_�a�#?�j�	o�D� ��!C7�*�3|}�J����Id͙���!5iѼ��v�&KW_��d���H�1��hb�Qw����P�!�
u(���KOA�O��b������}��Hbu��<���}\�:�Qr@j&!�����A�+l�� �g2"�t�Aiv�6μ-+o�z��*�*#-�X����u'8��E�,�d/�@�w�k��*�^u��~�jV�{������΄}�ۧ��]9�󗺀vՀt�>yԘF""G�x��CL-��Ы�Q��ɫ*Ŀ�����٘/�<����QVw�2�$�{p!
*�?���Z�
�4��7�o ;?���R��0� �YQ�&=�	K-<ķ��š#��1�`� 0�zhWwh�:s��~cd����U���\�S|��(q��ʖ��i_�-�7u�x�3���� &�]E��[PL�c��3jn��)�Υ�k?8�ƃu���3�f��f�X��Vd	t/<�~ĉ5��B��	@��3��Z���"��>���ω��R��VyG��S�3�c(J�=?RKZ�Ch�Ą<6_���W���
D$��p�����F$]��tSJS�/VK�9#�/��8��)x�cXyB`) w�����C���J���~=�u�;�C�.B�h�9�en_�¯+��G>������h�����j�J�&ߨUC����TD��T�� +#���#��<&8��\m�L�=�Uا@{I�^Ӡ�y���	K|6}�Z�1/0j�Kl�_��'�_uW���kq������j0��Y&c�Q<�FAn��F�h�Gw���;}��ս1j"�,�r�n���#<�F�(L�k�yxR��b��d���*>�̻�AE(t;���O0�"6/��[���DS�6h�dH�q=mk��R2����ʤL�婼�6j�QZ��)ȳ��x�L����5����l_f�al����b�)mu]��}��-�yh�7��Ubk~�{�H�4r���������o�����o��-�%��@��y��7����8��Iz�.(6J���s�s#��k�*Aw�9X��:����t�)^�ĉϳ�tJ!����h\���״�͵���4����`:���O ?�Gf�K�y�Ъ�3��o/ɸ�:
<z�t���
�m��Ά9�6�<��K����M-( �� ��
o+#	Q��UiY�V-����P�7^�Zf�H=~�U�sg�T�&�����B����$����M0M��5X���0-�� c;-R��$��-�Qp����G�vE�)�p8A��B{U�{�	ks�8ά^�R��Vx=����S�Tktkh ���'@��̑�h��#��΢ɻĽ������C�����J��W8?b��rV�8}��ˑ��\tR�뤊�e�����hj=r7���&k�#��v��;�@��̣�yJ�%iZo��;<�+��*�l�>�͉3��B�#�MN�%�����c���Clg ��`v�0��С1⡭�c]��'��/��'�b'���jf����-���N�����l��SP-5,�xw�'.��Y��A�� ���~8		��ԕ��<7�[��c�uq�RV�#��N�Z��k�qs_z��?�- ���x�%:��{k�w1�/z{w�/r19G��/�b�(���t����Wk�b3rjy�x�^k�{�*��t��ֹ��
g^ "�gD:����rX��K����(^�cꥤ=����uJ�e���%@a�
�>9š�P)��x��n�l�[Lb�1�N���۝�p��a����̸W���G�f����mx���V�1�i�����opy�.ùA0����)r�Zf�q��є_R��ű�r��������K��\s��`���B�掦*��ΐ�|�X���{z݅�9B�ߏ��vRC���f�$��b�hRcǉ�U^l3n�*��R'U����F�5;A��ԷU^��FU�`�YVQp$�)�� ,Q��A��-E|���V�Zc�5�'6�8�p�~ʚ"L�j���2�,cTJ��W�P*"#]�zZ'�[�n�1]�\�d��m��62�O��%�̖��H��r���_���Ǖ�l�f��'���Y���C���ۿHF����	Tϖ>I@����?�q���`t��5a4�� [{tE�]-�r�@M�N��|�5g�~i�\Jum��OaXs�� �Uitk����UE ���3W���+�{Ͽ�|U�p�7��(S�xѠ����Y�����AzAPkJ��b������k����ja]AY_P&�l�C��FQ���#��wC���i�3��H`
v.4z h`���F�f�'�G��[��:bV7���)��4gs�t'�F��ެuTD��ϻu�?��a�,�*d:��kԩ�+f�����(����[��bU�M#���K�y1L�����J�q�!� �+�&�!���Ǣ�}r�s{O��w����s����]���p��z����\��-��k��3�ӓy��}��рߝ���\M�*�����5K�Z{)����(��63���̭��j�<�Z�O�b�=��o8g�[~oBh�)��� .<�u�P��)J��v���T��ڑc��̮��?\��Hb�~!kWglK2ӵ!اE�TL6����@N[eb~����ԙ�v�4�8R�;�P�	B���L�g7�ȗ?�_���#a��B���8qsW���s?Q~Q�Vk��3`�*��!�/m��Q����÷��|��/.�IV蚨G��������}!3Ҥ���
�Á��up�G$�EJxJ�+&���_\d��������uI�g�������uC�8}/���yO����n�`�`�(r��~6�W���צ���t���K�S�fL�����j_���_�D>_�m�ȑ��l7��ry{E��
G!�[�~���#�#�:x�Fݳ�i@|�����
�|��뻜������aɑH�������m���̰k����JE ����3#�t�D� w���Q��<�ZRq����jw��ya��l�u����r�9$P�ٲH�z�{��^?�n����j)�E>	�t�ש��йU~hcp(F4Ί��}�(W6MWF���B��}!�����;ݜg�z�J�f&	�@H9!�j��c_0�[�Co�9!��p��]�56[!����mF���̅�onl�����x3�g��W���Ш	�=��ڜ����Sy/�sK��\������B�l+����T�M�[�W�O�&`m��B���҂p�ӳ�%��� BI��5Pzg��W�����5�Q2�91� C*;��)�h��-�h��)G��W��H��^Kn�P� 7��A��U���L'3Ҹ �bl綦U����j_�����?��/pR_�
�����l����v��d�Nh��[!��ͧU�����b����n�k1���Ʃp��͕G��2�����1��)�Ҥ�:ML[*'i�m�ރ�.x�4-Ru���U�F��������v>�*gW������S�1��쀓=�?U���rf;t����l���I���A5���S^PI"ƜRV���,��'��K�Z�P�?�����;d�p�S'8b�H��SW!���uX3�{o��%e`��*�Jܧ�>/���\-�a��J�i��[�>�����Y��r5*�>��֮��}%�A9�zR��`u/E���|}�n� �.vq�l����)��f$C5X����Lˬ���$��HJ7Q�	P�MX��v��ѽH��r�`�kET�7�?���r9c)rWL��z������Xʷw�M�ݝܠک�̳�tEJ�rOd�LZM�2����y�I,��u�I~,�u&BG���?@�-�M�v��wi}�l�i�a~t����ozC��K����������~���$��2�ڑRoǷ/�8t���\N�X^����TC���K�i�8v�EI��5hm�*�:�d�to����"�z�;��@���M���~q��b[]B�e�5�qD��}����������e��P^�=�X)��ӫ�=���r��r��W�[ k�i���Od� ztJ|Ѳ�γ/�1B�I3o�]�[���t�y�������X)�K)�!��tw�j�S1�U�C�r�1$6�m�L�`ab\z��Z��r���N�]?R�g���~0	�.(8�=�h.K�e���{�C)��{O��^�����_Q)%��u�o����v��O9f�+p�FH5^c��1q�{���z�r�'ŉ�e�V\c.3������J�f���eNq�8$^a$��t��\'���-	��Ў�G����]���X%)�X�C�xY��e6=�Zk��e�MK ���⦈��0s�/܃�>��,������Jj�\��:��&PJ5��+`c�u"��USݻ��{���@l�"�%��M����'0��e�q>'���� :���	�- �o�P�CdSw�:�<�s[,p���	f0%" �����"Kt2��DQpG��p�`��F:����Spn]�8��%%#�F:�Ƴ
a��s����iW��\�ȊU��Eꘃ�)d0W�|��Yu�F�~x��BS�@�oJ�|A�vڥa�	�j ߃q�_�k��ċ�U"Q�0���hM��x�^]��~=ی��:�g�~�5.�=�۩��A�x���'��P�k���O��U��C����7_P'�������n�Y��K��Ja�a�ws�r)l�q2�g��!s�n��B�^�����l��C���Zlb��*)G�9(PO�oΫ-Ro���V�5��8W�85=s�-�*W�Jl?�_�a>��s��dz��$s�/,u����z�C2����'/
_��i�Hf.��6+���ӠVm�t)�X�8H0���V(��̡��L�~�ݸ�*�Ϝ��q��}�sj�s ��bs�C����!�%����[��I�im��s�}s���Ҷ/P瑬�	������� ԿA�	�?d;����	p ��&Yp����;Y=���W���PK���/�V�2�fK [(XȘ �6�8��z�v��_�x��&��b��͖ʂ�����
*';p��1���L�Љ4�V�j�,�5�$a|Vz��o�%D�'�l0b ����IC61�L���d�8f�
L�ک=@a��8���_��M��5:qZW��o��1�Ǻ7}�b�P^�(}?Р��7�<��@�e��o� h�r�])�w�c�2~R��3�͊6���?3O��ދ����]d#ʱ���D��@�O)+"1��><7W�U��
6J��}�׶M'�[cZD� )���]���'�x��.��P�� ��Z�BSzr,d锿*�9�y�pOi���=��r�GD���:uU�-m_�4gb�x���Ӱ��k�Ne����9��J�4,�$W-�f|��e�i���EP8ҳ[S�7su��τGQU>2�֢v���;W��,�8#EW���}�Y��է⭽�U�r=�ڷ�^��T�Bɱ�O{vS�ݦ�Jb�Qc��K��~��
p:v�5�x>�e)T��lF{�#���ב�"U;�A]O=�E�w�^�H��~�F�`��8���%)*`�d�.�6,��NƔ�"Z�9�8>b ����K�B�!
��4b�]�8'�ŕ��̨�"ώ��.��.�w�U�l��(B�Zh����,�ѭo��>��ބb~�y�FY���hs�`�^����^��M�p_(�+�\Ŕ������An�g��;`=�D`��O���Q��|�Rw�h��-9;b�T�J���W���!��؉L��U|���>A��	�V��1�beZ�m��d���F"�8������<Tamϡ����!>ͷl�C� p�%�X�8Z�J*=F�s�� Wzy�9iza@ڥ �T7���h�-�S��9	C��cW1ݫY]���^B�Y� a���~-��(l0g���p�M-�';p��8=&�ӈP1���\<���焯l����Apc �/ �M��7�ƌy/��736�t��B�lɞ8�@ÌB�}����x�K�0��I/��v�\[�3L ���s�Z��"l�g[Ŷs}2�o�W�)Bt����,�)
z��ْ��!����k�t>��~�����e���Rc�6=�l
m`�ָ
�������O>��9���F�rT̕6��Wb
x�s�J@��aIH���~x�$���i�H�%W&W�,������J&8��k;,K@��i�
��C�/�C���ᥥ¿\��LTU��G/�`�e®���6h�p��SG��N`,N�_k*�h�<���+��(�t�-e:�X�2,˭��,�c��_x$�����Z�(��'@�Ä��}�W�,J���X{ŭc��`$�Wy<�������T��lK:��y����^�ǹ����\2g����m����%��O!���U�-Z)�ekq�/(�"�L'�'����'��.����7�}�t�x����'m'�7��)��6ٔ��۫(�<$n�j6Z%}u�o�](�����J�T�~V_���x���n�[�{*��L��Õ �|���i](�7���׆�վ آ��6�ā�m���hA��&w��9k�47�P�g�!�2��Q`{q�F֒�}���{�ki���d�*�uƑ=�cq�� o~�ۣd�2��>�T$;i���@��z]����?�_1�1ɞ���C�d���G3��|�\��*t?	��/���ՙ��U**&ٸ6�VO�%+�ݼ���m���d�ɂ�I�8.��pg�H=�؜�9�|]�h#[M|/�]��3<����L���,�I+��q)���.!����;��\r&��6_O��ukI`!�v�V�5��E���S�"��+H�R���ޢ���[[f	T�C��L̨�?oJ�i�)6%ep����B:��dD5|z��i�#�巖+��ʵ��8Q�Q��$>
��O��F�K(�������|�O���7*�v`��v�"}�ID).��� �!#Uj�|I�^�f��) :�˙��j�ZGYE�,�o0�����S�����o)��2�{�$U=i��~��OS
SEؘ��;�[\
����s0�ϒ7�'b�yJ��x{_jMӖ|��b;'DT1��K��u*�L2��>C�XEJ#�9�^��_�]���;�D����,��3~+^@�*]��������s�+��o\8(JTC��=YP��<0���^�s�JE�z��OO&����p���R��r�@��zMl����~��B�����������e�)���ֽ,@Uݛ��A8���/M�&�C�s���7Z��.ؑH^E�93��r�n ۋ*�YK��2Q���>�fgq5�Ѵ6'D�s6(�Qk��g�<ϛ�x��ԎF�m���:Jb����f�$I8�1�0\�r�$P�OZR�r�OM�\B���Yk->��Օ7̈́�r�ܪD=����gt��uV�W����y�su��v8sj)��T�{T���,�B�Hy���4iJ�t��1���>�������8�Z�rĢ6¡�͎���Qj����a[�2�`�]�����8�e(B3�I��| H�a�1�Wt͹��F��=�����R�����9!}x�;:g�t]�R�0f��͢l�A��M�O7څcK��f�bO�,��q�~��]��)�pI��������*G$y}��ӝ�	��q�_�u��M�����������W+"r.�c�k���΀/���S��͓Q�y�!�ѽ()q���v��A�d�S�jp=61C���:�՛�� ��p��;���O���z&��8L�3-m�{5���ZX�V�3�1�Q�VE)��e�%�k���34t�*�ժ��a
�t	�:x�u��<Y����jzg+�+��]�\�j�qߩA̜x��^r^���(9�3�h�t��h<��M�!uo̴�F����_��BK�Z�w�:ю8��݆x���Ǌ27V�� R��W���0���Uu��S�6"}p����)��z8��#ȩ\vX�۟�u*\˱�|.pTل�W�Z�8fSR|0*=��&�^�������[|;��[�(0��E�a����S���|؛�K��9��缣��X�/2��r�ե?�F.5$��h��"�X�B56&���l�ut	���~o�f>dZ[�+��[�j	ˬŻ�u����"w�|��mяM�*��:xGk�o
����U,@o���oj)��n�� �
��G3G�e�vjah5C�[Y[{���^��L�M��`�Y�UK���ɲ�`W3�s-�V�]Qܻ�����T�ZXȿ������!�%e�4�m�
���C�����G���9��'l�%}U��R�֡���2)�O�/k�>�.��ă>�΢�V��V��#b۸��7T��N���b�v������#D�v�;0���8d!��;�++�v�X_��m1w|.}���g��2�R����g�yش�ê4��C��:l�	 n�.W#��5�7S a���}�r��[�h��-�bþ�'ժ�kN\\vXM����H����,{�T���}�o-S�]�c�,�̏�4��[\�9���u�NV�H�ȅ���̵"������u<7���ђ靖��jz_��A�fT+�u��x��%R/#N͂+>���H9z�=�&JN�/�������W&P^ar�Ȣ��#] �ު�w�~�Wx��LT��Fθ�2o�o�J[�����>e�wjn'�Yjbs�$@��8>���W+!?6��؋·�ʐa|�LB�a5{^���Їi`�N��b��^JBڌ��L�B��I�'�{�R8�35k�)Y�g1�K�c���BU�GO'��K+�Go'4JATL���� `p�⁳'n��x�U
]�4��:6�I�v}�f��������_tj�)�Rʣ/:M>�pv S�Nd�'�N/c�<kJ�Y ?�*�{L�S�^s�݄�@=�6�����c!6�<�Y)���0ݦ�l(FkI{Ŧq�5�BMq/��f3����+���ð�QJ<K�j�$�)	4�S�z�Y&�t��A]��UC�V��Dԭ/a콯��c����������8>�k��q��0��-���0c�i[��4�?��GU���E&�^���:��cG�_��/�ԥ3�Yدk]P����B���S�[jF���2}�zezQ�cݟJ'��wf���!U�a#BT0��U�weB�sQ�s��'���01�-CRg�5kpՌ�~������UA7��[I�#)Ȭ����G)�������'�Ĕ��q|��X�{۝�2U��^���鰨�${fW��Hu����L-Ǆ1kz�����0�HR{��[����d�7}��0
8�����-�갑Rx}k�V�QPĕ���y�n��yO��E-C��B� %�=�H6h�,l�C����E�^y���&D�ͅ��E��Ż���F�:ב�@<C&qB&$X�G����K)bH&�}�"��q�'L��[���Ͷv�A��u��7��;��?
�Z^i�
�`$'��T�f>������@z���h(�����2����P�w��160.��c��]?m=�%��ւf;#^����r3����Ρ��dpΓώ�h�}���S��s��:l忶��$�4��#J��P<�Ct�ݛ���t}����q�qU!�v���g�Q<�g(��F���O�zJS�3�i��l�s�J:/~�煓�:�t��W��V1b|��\���[w� toa�����wM$$RaB\vGo��B�פ��_	�w�Vޮ]	\��&�Ξ��p���4�J�p��	9|ĬE="�þ
��Ē�?|g����vc+���m[\ �E�o��e!����g*%���
�*��ΕX����dJ����� `�n�`1L@c�I���lӼ�\�MG���}V���:r���+ۄ��p$}�e����v|����|z�3��M����bW�5�Bb[J:+�������J�.�K�PE��!�V�CP!��l�#YA�M����@����Wr��}�@�mE�DK�q�ʼ�������S��:�D��M[%'0�{N	w�p1�Y�Xz��Ҧrj�0r=S�B��'���9Eo:3����Ƶ�	���例�F?t�AZ�� C���X�.�PWIN�}�y4D{�`�7n�rہ��N�\	�nQ�+8}ÿL�k(�k1��?�<H^LP�鷲5T�nd�~d��:7�G�	]��������8k
��P,�.3�"	�;�$���n��<�&�B4[��է	���2;��P���K����`�n82Y�g���6s��cְl�-��#���+���Qyc�\ЅO.H�Ĭs���Z��!��oҷx���y[��F�q�F�L-a�� �)N1A�����FqE�i=}Ŋ�~�sp��)i�}�9��	W�m�0�X����Ct@���õx��2# �L!�#�K*�D?B�����c9���@a�����J�6Ei�R�m�rD�'�Ҵ�ǚ�qG�,,z��	�V��`���_����ɘ��8�z�=<aB[��e�YBr�M;E{b����%���Q�m�	�ȗ�O��d�- �ҚN=����s��)	H����L`��Z!��	rP4�*;�[3������e�2�3�?XU�}w�3'{ξ�i2'no;�yB��J'��}��{O�CX!�@����Wj3��VFf��ZhO��h�GH�Y�rۧ]�v���X`pu�M$d��W_��0��(,z�7cquiP9�gk���(9IKK;9OB�����Ma�I��<�tӦ��Em��*��~Cql`DIzO�����^�;�{Utѵ���3I�ðRd�i��ȭ!�s��2�*���/�[q�K ��Z�rm�˶�����r��~���
�D%�����f"��:��,��c�/](����?0M�okI�Y��S,a����B��r���؝�X㒒����]��iCQ�T�$��y���>}/�&���q�˻�9�����7i�6�d�ׇ�_���K�Uq?=Bw�E|��RC�&8]����(c8�^z����}U�M�j���Z���ѕ���]D��4�i^q�l ?�%ۻ����Mdr{/o����\�C(õtM���.ȱ/�׸��p�ń	D��!p�I��/���7�^��=�u���2�L��)'����YK�
��N�8�3���X߅�0���+�;��-���:
��8�.A�@ɗ���8�T�+��֘F��\,���)�:ƞ�����7*�Vu/i�v��k(��0���C�4��߇��W��D�8M������
��:��<�m����Qj�KU�������G���{���>�٨�rǻ�zٮ洛A�t˯�Na�ݽ�A't� ��6WKa�L�����&��]�����"�lX�;��r�sT��|̺��*v=��6B5W���4)�	H�1 ��&ɔ{�=iM�{������x�y�7e��s9��k��(��G����3��zi�-���p�	����g ��19�j>����Tɾ��:��k���7�Q�~��r��d{�
攻݊��1wĬW����~��Ԉ�X��5�cxkپ��4����aW�h���n|��h��_��[8 ��T����+�!���W�W����ln��Ea{�3h� Ǎ>�rs������N%ty�Jj �^��K�-4�+�ӆ���ٛ"��!�dH���fo�+(Y��lu�����|��/�ݡŀ�����C�ZL'&j����]���lG���`��3����o|�����p�����m�gOU3!�������je5m~v�\�D{�v�G$�%�x����R�<_�i95��уc1����~�&��]�X���RZ2��l^�@ʔ��-�#B�>�4��N9u=&��>���� �����[B��؟���|�r��}�RE�����}*c�������uFi�DV��ei[}\�2MƋA�O�j&'�a�֡j�w9!bh�8��=(��+S�
�B�i@Q��ng���AB�/�# ���Wi?�48,�bVW�\�H�౰���SC���@��[�A�j��a����N�,������l5�y�U�[��2��}0rP��6���T�
�ro� �
���[��1��+���AvJV���T�/K����a�-9 ���v���/?�[aW�Y%Gp׋�c[��^\fx�W������ݟ�"�k�Ӊ��P-Ld>Y�c�\%�U���3��n�gh#$ �G/]��ᰟ�}��K�J���p��18q��hlHf�����*I���G�kx�� �K_��)4q���oĲu���1E.����au%������I��C7�"J�,w�Ygc��y3湬���.o~���F��a'wg��vk,�.H5��X����i������@�h���^�:/J��Y�f��y��#��t����}�V�s�����$ۙ�A�'�L\��>���d���X�5Ò�V��h�߼�{�1?�@�7f3۹�G�=�Z�(t��ݛ�\�u�)s�{q��5����h����ن�M7�rRI?���{ܺ=��~l�s�=��}7v���K�}���[�8@�%�{CPlL+5)��qC%�T��Z9�X�g�/�Nߨ�gU-	��T/Isaѳ�)n*�h�� ��^ކW-�B/b��?�jͿJ/:�Pc�VҡѦM����'`f ?�G�ռ�ܶ�*��41�L�v��C�{wU���@�v�h �ӳN��9
W��#��\�_�4O��#*i�.Yj�<�v�{kxTo:�`���&�^�k��95p�c��tD؅�ᣔ�;v�)r?pv��so�qj��Ʊ����Q��p4֬��\��â�l��3Ks�J�swM>`�x�IM�?�l"�� ��8B���tF�(J���)�b�TL\��&�❰/��KJQ�=���=�4�SX#{Ҡ)�/�R��X�S��tˌ�8���E�QQ�<��M�]�CN�;�X���5?�V���:���Tʪ�U�|Y�cR���+yvi���w�����2�)�yS��:Y	��6 gv�����;�[}֑�눋��PZ���&��p���Ү�_g��,x�M^OY�z��Sb�^P�ݫ�~��Uڞ*^}t[Vw[[ 
���^�jzi�m�'���_HO��BvY'b.0\�������'�7
�~���p��wče��������?nQɞ�t����w�|'>u��*[9�}K+}p��)?��K�67_}�]��M�BS%ْ!��n��@�������.�zq��ac)'�I�C�n5_����v�~	b�8��Z��֭�e���&Qi���K���|�OV�$j\�a���4,�1/����V���^��p��Y*�v{��i��Wn{�h���V�dpX}Fس�WI��m܊北��(+3°�Fs�*hU�H�� �E1�j�o�'d1oW�a���d��0Lj?���/ʻ1�hl%�x�������Aa'�~��H��0�@�X����Ћ%qQ_M�K4��T:_x�"��]
;�޾ֽj1z۴��ch�Jx��bQ6!߇�J�=�4uhܖ��thE^�5�j׽�]��__�W���B��ܴ��樬sbFrA
2`D��uz�����
�Z/�s���7���"�*_C�>���ـB���}B� N,��Ut�͠h���t6u�f_\xU������-�(n�Q�_����͡Zѷ�$s���ү�ۣ��`�'P��X$'/"2�Kzk$��HY��+�)p=��&������q�6�����X�R�n�f7�3%�4�N1�ڨ�6��	vw2�ࠒVӭ����8*�I��\�\p�l6iMxЧ�v/���*��M�Y��1��+��mW�[H���g�@߶��Ɂ�V���kE��C�����I"]�6�	�ڛ/H-���-Zi�sj�K��t[����H5@��H�~%9`ދ:�s$)�Ƕ2�D�>NH�X�xB���纊� =�p�þ����d:��K�Б:�N�tR�����lcF�dA����SӫA�{A�D[��_	�$PV>чI�T�Rs�QB�;(�\䡅����)��!!�|h��z���p��L	!a0��*g�i��24Di��@-%z�Uu���=����3�{ɻ����W�c�	��
}^Y}f�o�9MlqM��.W@�������M2�=!����$��	KKYOt ����ԍ�JN�%[0E��	�pY�����V����ϑ����Z�ͬk����ȓ�$�u������V�N�{�@��6�	a�Wo?�ͩ��[�AӔӜ��YcL�(�b�e�w�%d��19�D9y=b�씢��A;�;҃�)��<k��<����-E����xc%Znǲq�$�wo���%���gŲ��\�ۣ{�>?R��G�����U�ҍ�U��'���o���Pn�����s���ܟ"��H��<�o�}'Eb닍��O'�xc{V,`5���jó�t�{��g���
��JH�)���t�Lj��F��p�Z�������jֲwL�u>�Is�#+�5!�V�$��˘��)�w���}�'�
�L�����#mo{(��"zFg�2˿T�.�ZH��H
��D�pt�Jӟ�Erل�V{�r8��F ��$'+(�T�q�O��qB�X&������I־U��#�q�^�����E�/�%F���qU#�E�Q�:��a�H�aԱ{4��ot��֗Q;�u�<ui���z��=�E��<���D0������VaxK�?:�1|���3��٥�W�����L~����Q���J����L��J�E�\�z7�o��=L���j�O���6�x.�۫�zP�!g�c�M��ˢ���mg���ڵ�"j��t�lhV:�~2�ұ�����t��9���Էz-}=�"2aL��70�Uh*G}�0��a�	Vr��WJb9V�����m������zؐ9x����e!Ԁ(?������}� ?=k�A��Pw>b�JrS���K�c�Ѥ^T�2
��8a�L��,��L�Ħf��W�v�W�RҖ'.��V S�>�;_�����e�}�[�_��i�43��r��Cͭ|FL@5)��/0��bzK��ĜO��ڍ�łV-vG�`���つ�7���!y�e�W�S+��ww�ɞ���lz+��Pd��_��EH��fr��
2��]�Y֧	��3�ߑ֦y��x�#��/���Y��Ѻƺ�N�k��'Y�'��A"-����,;j>#uv�`h3�?!��E��L�w�,ʨh����a�[_�TC`"����Zg����_�J�{A��_ʐ���M�Վ��S���pr&�@��"���l!,̻O��p�/�33�i���K�'�n7Δj~5V�
����0�K�p4҄�!��[H��u,g�G'/�J�H��<���g�Y�?� �>?�%i��)8�-,�5�ut|�N�J���.�Z�u�X�:B�حF�A�+����l�L�R��*���[�FG�2nI����@��u,?�%A�~�x�^��B�&�>���-��x�(P�z��P��h�D�K٧g�*8���dzv�`1��EX@0X�t(rϾ��1��$���`B�T�8PV0�D�w����H�d�>Rt��Ѣ��\E�_�+�+׵{Q��R@a]��:��q#���:s?໋�����*��̱��|�܂!bN��gTToٿl�]��S�#�Y,\<���Ek�z�暠
Nؕ����x8l@-��U�*���t�W�f�H-�z,Ȑvl L_��`=��\�� vZ׏�H���<�Cy�5�LJRY�@o4]�fm�W$�$
j����y��6O���\e�e-A��8W�V�8�AX�ͦ�r$�疭�;��~j�h��7��[IOX���		���j!ʺ�?��jQ<F�-F
��=M��E)-������ԡT��lc##�vo����q}Ƿ 	��6�bB!�t�u��.����TP�G����$�$oa^LK:4h����	�+S�H�B1SX1a�����1�Ƴ��r�ک��c=^��K����$���/�Í!��B��TY?�H����0�gzS��������Qr"��}���ގ8��S8��?�p�~N����x(?Ï���94����Y�Rs�����2�%]a�m�b���x��S���jA�c_��)j�j5��[;q9˅a�]ڿڗ�����&1��?O{Z���2ʫ��ǻ��B�}��8PKO�`�e�[��Sol�O���<s�����/�ꄈD,㮾�ks�$�6��
K�A0��Ï&L�EF����8�B��[��h"�f⻻^ؒ��?ЙX�lMs+� 
R��S�ʁ]S���6���y,�@����uj���+#�š���� �(��Ą�*`;���4|Ksd{�kL:������M�"�n>�y��WZW�>֤X�Wf�>ޗ�J ⩗5�,,#@����u̾8e��Ͳ�$C����z�:� T螜Z����8�s��Y4��-��,�(�
��{�������4L9;U
������΀�OqUM<�f���_5L'�0[ͬ��(�S?)�ww���g�5�u�/6��~��~6��}}:�;�n��^Zk_�$i���1s�Lz]��X�8��9��ƴ��q�h۔�^إە��ڭ�X�PHz5+�i��M}Ñ�P�4;��qn��\.���&�!�Ļ����5�c
�a"�<񎊐�яI��"����>\[�0�*[:.L��@.^��n#����V��ܻCA"�X�:�ېĕ5�*{��;��u�ե�L���+��|�Mߞ�y D�{�s������ϑշ�YIH�i�G0]<.�k؀U� Wa��f���4L�aD�l�!LLgk��U�)U#BP?�y�-���4�"N�� �����iH����� ��z��K���öNZ�TO�f���x��S���t�[��>�-^|�Ŋ�L�WF�Bc�]�����B��iK��];��"ɟ�_eHLh�	~h���_��r^���Z���=�.��7({��JY_{��%?��}�HI��&C�ϤyX�F}'i8>^�#�U�"O�y7y<�q�Ai�V!����"_� �^QJh��=�˶�JP���ԪXԻU+G���yc�.s	��)Tn���AX�K��w|�}c�܋|��O�⍯,�&ONP�C��;}*�·����w�b5Y��V֧�ٷ��#
-�����"�%*}�	��w쿁Z�͘2hvc�W���B��Wf���&[<6��,3SE?�ϐ���[�0KÖdp��'��w%��F�$�%+������#u�@-�毋�K#����n��8=�aѵG�zB�?�*ݣ��8�s_�i�XW?6v1�͠?&R�� ��r�U���L�J�`+~*Ȩ
:>�<��|ت�b��%92�b��ye� ~��MǸ�
�Np.\KL_�q&3EWꟗ�&�v���D�O��A�Q_7�dcez�wP��w�"��V����^�H���B|6��ɚ���.
t��Sz6>T���Nd}aa_ܮ����� ]4u ���Sw&\kP��:I�l)9p�[e}����8�����ԥ����R5Y����r�hh�)�7 �0����FDx��_S�A#%.�p���#*)�͑o�-;Ы$����tx���I������8_�7 �;�����bq�2Ӗd-0c��F��B���!{��j�D�Z�7����7��:;������g�:o߼šޟ|�^��<g>����v��ڟ����[�8������3��K�W'3���\�|�؃�Eh^�2g��E�Z���c�!u���[4���*� �g!'qC�it����4Uͤi�n��L��R���r�?�m��M/��O�zڕ`_|�����]�o���`G��:��y�_Ɓ���_\�h�C�_zr���K)��e�3d)��bJ��ZK���ne�G4{�
��pNَ"% ���?��e��p^��UJ��떈����v�26�%�� ��u1R������&�࡜�R�ϸ�U#1���ps�x��"�����Fb�� �
����Ɛ�_R�����	�;j�i�%�e��^��֝����&��:���v�6?u��Ahe��/~g쁓�W׏Sm�3"
�.�8�`<B8ppz�>���#�����sy�Ka�����+��%��� h�*;�'ru��Р9L>Hg�<�LJ��vi�Z�
�-:��jƳ0���v�ty�[�TE<�l#��#�}Y���(ު�f�ԩZ�1���ǈ��dPZ��|-4�ស-���0�V�Gk�U^%B������;��*3�b��[S^�A��;	�x;���!7�O51�+߻	B٬�~H	�sld�gAd8t%Ά]~�c;����4˟*jF�cɫma�]dq�n*דW���A��� �'�ڹ���N-1=T�0��w�u=�ܢ'�X
�fMR�>�JaUu��{WG,�6谞�,�*�E7�$Y�z�n��i���[N�K�����7�!����eA���X��*C�]�}������!/���8�»f��a]"Wgq#3Sд?�l�z�����k&���XՖ�J]cVs�'ʉ�,��B�[v}��b��&�%H���B��S9�����[���N�����ѵ�0�P=�G���Ui��{�l.-�:��ƺ]@����n��w���+C7Amo+���+��Z���4�M�P�`^��#��e�2f�G,���2y�6x�r?(���Q*���R������ᖜ��/W�21��z�,���K��͈��K�]�k��t�zc`�T����P_�5��oi0�@	�L�~�I��Jp���@� Ξ���'��R��t��B�d��F�2�;O��4�!�E6��Wߛ@�� ���J�8./3���N�6N���Y�a@�ۡ���r�6�`Ma/~���긯�e���Vy���XJ�ބ�ֻ;���3t�p{�/,sM9~] U���tZPs&[1h�=|�M��N)
�b��`�p�ˈz�Xh;��6Xؾ���!�5�)T�-a�j�/uX�l���҉��@'��ZL��hDWBTl�nSH�\�W7A��������h$�E�~��,����C( F�#�ԥ�7�c����A�	��*N��;O����%�X����=v��J�x�Q��	�o-�*���w��wv�� E�(Cz��maǛ����u�Aݮ������n�Ԯ�B�c��E)W�l��sgC��&��WטD�==�$���������f�L�߷#�/�:�.���n��ş-A~.�\,��J�,4,��:p���a6Z`<ql�%R�o��PiR��]8V'c�L��`cmY�J ��ExUy��@�t�|�Zܽ6%�gx,lW��]���W��s������x��]�7]��g���)L`8��E1X+_j;Lעȫ��|���s(��Z�q9Z�c�AC�C�X��3�+o��D��Rm�`hjia5��Y΂��!�'�=X{_��ުX��/L��q�q���ב��W�e�)��L0��U����3�\&>x�EAb"��K�a��.2̑���2��d�Sq�Z���XA���� ��q��O����q�h��TG����|HQk��"h��O�"����7M]\����*�����2�(�"Y��j4mؤ~���l=��5@]�uO�X}r;����¨��m|8����WQ�Uc�
g�	�{�YZ�Afڍ�[S3�F���p䠏c���\/����B{?��\��fZ����x����Ѿ	�&%��ˬ�جI��/�Ąw��u�#bU���部n7A/��5Y��v�Ibg{�Z�����m�Pu%";+���=s�#l:��Ycy�_L@e��]�E�A*m� j�GV?��C-������U�uS<� U��\!��n�Bc�M=��g��B�=ű��~ɼ�w!��b��#zD,�n���d�QZ���n��%��6�?���J��|��_��xR�sr��{�<����WK����G��J�=$�
$�=F�u�P�|�	N�����I8Kӹ�ՕD�}!R%'��$DX��/�����C��'/��4=�z��Kq��|
�-�g_�6l�s���N�-�RIn���O�՗��}ɍOK�isGj��K�V�SR�ˡk����p�ԑ(~%�`�3:��74|w�N2&��?�g�MI�F�҃�58S����k���HXD�
{\=�h�����?��z E����Xşp�h�Zn��(���߮��HT�"����`ey>��k�d�6��A�Qze���/��ThWzbZ�"�����0>�ϊ
��6i�s�ZN*r��,�4���P��(Q4UT�E�eX�)b�w�oIr!�5�>��\X�lk,֡�8"PM��SqTz��J<Dh1������J�}�Q����w]b6m��j��!�s�x/��f1�۬.�ǩ�;0�%\f2s���ᐙ�O�D��pf�Ѣ1�H�C<�.ש���׮s$�m�Wi?�����j~p	-�=�M�����Δ��.'�\ٻ���_0ń$�����O���#W�Q#9���Լ�^D�%E�՗R�	/��Z��f�6�ߟY Ƈ;g@�_��ߺq��Q{@�ҽj�Q���Y��.ի}�:��r��"�L}������("pj�@�Gz���,�{��N����0�3��%X���i�*��ӵ+�ߔ�@�/�x��1�T��;�ղ]$�N#��N#G}�0Z�/��p,���H�E�9T�i�'С��I�fo�ş�^�<1G:�,qh���P�c�
#�u:8��RS`�e-�uy["�䲻u&T�$r�1׽D���݅F�Tq9j���E2�a:�ʿ禋�$E��K<{D�=9c�I����Z�$J#P�7-�*�-;/:�ٔ�EW�䲁���7>���x�Z�tD���8\�H�y���"U��׫/��>8�V�$���@��jq��ծϩ��~7��e�����*u��:� 9ݍ���#�%oE@�e�p}�2#�I�B}����K~��ξ��� _ف��r|���ro�$P�\���)�[��z�c7#*��uϻN������f�8m�og�ѴS�r= ��b� �Հ������K�p��XV� �U�̃jkuF���5���h5&�|�u.�4T�=+���G6����Q�4��v���p���a:�Z��oTh�(7�I0|io����	�VF��o�r���W�'��ғ�@M�q ��e�&�n�;ƶȬ-sc�'B�J�����0��uW�����c慔�q���k���r[������v*�L�-a���K���|�wC�T� )a>��Nx׵ `�x����!���]�O޳�r%�+��d4t+��[{r�EGi��XC���N;�q;>D���s�S��f����,|2���8�I]9~0�H#`��yg�9ZH��D�Si��lCo/�Wr���������`O����~Us���
3�}Y�2�#�m�S ��� �3�YS�!ӫ�Ng�00����
���`28٭f_a�z9���{h��3 i�'=�u}���g�
�8��N4-�S��2�ک| Wį%`�����y�_}?Sr ��72 �s2�4K>ˀ �2��v>��H�b��4̴>S'x�#b����&���a����|��W֦�pv!Wލ����(�R����z~��Qv�H���7��+����J7�	�[�US(�̟�}���+������"��ĥ0-��%�vh�MqNF��+�*6j��%|c~�f�☳�����q &j��s^��ܑ��6�a���ЙD3b덐l::�㽽=��ۡ����,�<��ֳ�B�b1 �6%�)�}���ʄd1��(��-���\" �ǱpE�	S�oc8�f�FLY;�Ĩ�������}L�D���Q�`Ֆ+��$���װ}��v���64�fb�f@�˷�-��j�!�Rm<X�o>�Y�ɩuSl��2W��������R�'��<2˘8�=n�ڭ��Ч��/:��ꔼ!h[d��S��\�J\q��c׋�A飛2D��y-P7�$+��B{q=�b�C����g�~����M�1����F)�K@�l���r�>����b7�+�\�mҒr x�_N=64�A�Z��8ݒ���f����](+���l�
2���#����$鳰(������߈6�h�l���ǒ����o�p��s�`n�@*��#'��W��=�����;k��|�j��J��V��Y@�A�$z+r��2d���;;���9���q}�1,\��GƢ���1s	�����	h��f�!;��Ռar�������m�܃��v=�B�}�΂l�fX��!>#�ѐʣZ}��k�рg:En�9�lJ5�d�,��Ȅv�m�1�/H�j/��%��o��� �f�B�aڿ�dݹ�,arr� E,N����P=��^��K���$�tџ���SA����Ћ���R�ں��:e��v��$Սm���Q[РӘ��Z��<��,ֈ���6e?�t�~F��[��iP^�M����G�B�=�6e2���-����5YS*��+�:�]��	&y>�3�VYߛ+	�@��
Qj����������q�G��ɽ����;��O�`g䦟���k�.d�gL썄t��d|����c�h̹�%���^�R3�I$�OǆQY쇴��X}��ЍF>�*@E�9�8�<�B���&*��bja���W2�0o��y�r�ҳ�1y�cXx;p䖃�`��$n��D���΋��2�Szti���C�>UnA����ߴ=`�d������M�ؙw��N�lA�̕�QN�6a�
�f�[<2	s�M@:6��$��o�G��)�@�x�x��l�&/�p&&��dB�����{�-'�,�|a%yȉ�/2�['���b���ҁ��`2�2T�لf�-�[��"Lz��r��)#,Lxx��ȃ�K�
k�@������1��������]�;�x���A>����m�j�sYX��r�_���T:���F<f�G|�/�Sh{T|u����{�=�/����>�4��P"r������+a�ޞ�K=��a�i�������Ls�ɷz�.N�Ly�'�4󈓿�	�wbSC��ñr���Ҭ#� d���PZ����1 ��M�hrr�9�F���Q7֦���˵`
f2r�[b�0xZ2�p���`�kY=�q8�͕j��S��&Nu!�����@ )����sB��+�??�I��G����W�Ob�&��_61�@U^.ȵx+ttB�L�b̘Y���c�E`�/��\r��i>+�X�F7���wR8�䯺�<&�:I�W6εtH9锕�+G�B-g��{��H�u.������\3��[�	�ɡ�/�XK5�>���cE��t��2�&,:�ܣ?w�V�ԏ�A��Y����x�$t����>�R�ZƗ�t���3(�	n&�tF!����V�w��v�9G��b��wfʢ@��^|v[Ԗ�≳�Z:�ˡV�
l:WYꁱ�D��$�L�����m���\eJ#K)�L>,;��/�t�J����DZ��r���ay40X�\e�sa�ΰ��
�l���h[��!�s/�n!sqz��wH�Z�d�C�5�U��?�Ӹh�����AA5%v��8u�1w����~a�hF�X���ݬm��3��c�Ǉul�;�^��)bτ����+�@>rRN�����߻��{�˄�V��sfӊ�b�Xw�����o������'�%�~������}AG�,��"6�g¦��$]�h�8�}~��l�`�����X�>��-z�9|:�3�+�o�.�3{������3�ӕ��Bn.l}��!�[�CԽ��J�2bn����P�9?!:�C$
��P�S��8�BK��Y"��ܴ��I���6D�z���F���C\��AܕH���(G��C��<7��y�~*�`a�32D�R�w$5�&�e!�)��7�!�q��d当��׊R{�mr��Z��f��4�^���q�
�����$�����>�UTp�C�ݭ&4]4Ӎ�}���TB������d�p:���gٶb�[N`D���1�N�d0��4�!�c8��~������t���Jg�q����l빊�I�������N6aŹ�s��2�\��Q^_XwC���=M�v��U (V�ئz%�6h�,��O�7�w�Z�2Syp'��1 �X����M��mg�D�4�O7|��-�#��)��ݛ7��\Y�}�2U��d�;L����~&aF�c�?�r�=2:�m�52�ʯ,9w0ަ5:�i�yDX�~.2�p�7���&� .Z�)~C�(<N�yuU�U�?�X���u��暕u�y5-'�������������7+�(b�3{��l�����&Գ)s�}g��^�5�b��1w���ԱzQ=�W|��O���nT0��x�����!@�RsX��?}�7��k������S?l5P��Y�� ��ѭ~�}˓�
�ό�����F�Ly��r�'0�ʐ�E>2�5�<�v�n^9H#�9_�R�6?�{�)%��%G3M%8/3�K���5T��:�����@Bɂ;*e������$PP	0Q���j����f=Q����,�T��j���;֘6,�k�Vn�^�h���"s=��)�x:�/��s�Lz	�,�[��)y ��fOgmn٨�صt50� �Wt�����u�Ä��	��{��^Fc��#9��t̅�̫�;���m0�N�f���9�uZ�+/�i�����y�N6�R�e?̧@����G��wl'd�z݀���C�E�1TE��I�9N���k ���V~R_؝	�i#�5�'QRIj8Z1�'�֥\p1-�kUYƅsC�]V�]�d��哦o��l��v��ɠ�u �����������!e�0SZ�M7�${D_��Ѩ�&ja$Qڨ��$u/�.-�4j!�������Ǔbj*:h�W50�����z�{>�0�0��Xi��T?�Ԉ��Y�%���>HDlx����`��`hmuO� C�.��~@�z���Y���<ds�jj9�/�=S�2��v�X��ԘZe�s���tc���� 7Y�[z} R:��6��>��״��+�o�V��~�{k���)a��qI-��k�[k)Δ�ވ�:8Jg� �����L���C�7C$�L�'m8Q:E��&I:;���/?�M��L��-���� ����sV���4AF��)�ٳ���ϢC��2�-�h	b�>�֒�xH���N)�/����� i�r:c/j0Z�e�;���e�ˌ�{�F�&D-�Ru9�8v���T%xF󙋕�d�F��r���w�<R��\��>���}�aA&<��R��
]���gD���B�Dչy�'����q��������|�Уb��H�}�\�x��C�����G�V{ӡ�o�- v4Nn���%[�	�ú-�;hv��������I`����$=?���?����q�Sg 0"�<��xD�%�����5�/���e]O5A|��G�D��9������G)�:��=v�2�,�;]�UA���b���������:�td��,��ڀ�����U8�k�cy.����+��L��4��@�o��)����Tl�Fzu�v�sM ��ɯV�B�yv: �l�ܺ�xN��� ?cE�@?�	�N�Uj&+,����'�+J�����T��W�lf�����7sP�d��^[eB����u'��g�3�6ˬ3�;XV�p�ct��V{��r�$��ي��\�]"��¢CR9�u)j��f��z]Π��T���o�1%Y�tm�9�f�B[�bG2�om[�V�_l�(���5yF�F�uF�����k�h	�x��v�|(�є ��A�gI�/}H�\Ŷ��z��/��oP���m"�I.�'�g����.���c��˾*Q��.��edF�o��[S��-Y1���ɭ�M�umd�Q'��j�-ߍ�b��=	��!v�dZ����6R����#jg}a�+on���i�o	��~n�+\t������Y�D��K�)��{XC��5����ǋ��F�J�R@�Zu��k	R�C���ہ9�an�w�>1G<y&����b��Ux����S~;S���D&��2��H�X>"Y�����	���5���ڽ��m=�(m������e���S�'yw��Ѹ.gm�:Lz��wj����t��_s�:��qH.��S~���w2HX�v��i���.G��|��:��q�M��gr'/�4�)*m�IC�'��<7�SRG��"oʢ�d7��jk��� uY���V�{Fg)���ui1|���~�`+v�'���-����Ȭ�Uɒ��Z�BȔԊ_��]${0,8RT'?�� 2���T��� 6�����3�A/5�3wb����|�Q��(F��G��Q7,�(���Ul�nW���J'�w����[Z%&TA' �i������EW .Z�Ie�d0�9�gc�� pfסw^}Xqt��-�k��U��[��<�y���)�*=]�@;�,*US4ǰֆ�^�ߙ�Rx�����HR���oQ6�e��jF
v�$��q���R�H�/�0Ɵ�O_y��$��*���vs��5�b1E\�K~������	�A�p��v0hE_q3���Q ��U�֘Ȁ��JgV�ʏg����'��p��I�J@D�]قtq��r<�r̡�@p<�͉�-� �J�a�9�wZW�^��rl��=��6T���Ycj��;e~M��9C���Q�����(\s�į�������BC/s(�eZ�[���2��)�u����/���d��R�ax;~�r�Ҝ�A��)j��τ�^utU���o�����kӚ�!JSnV�!&�� &�έ�<k1�u�`���u�dN��[���v��,��N�'e��2k%� �Ѥ�)��P��G�Ŭ�%(z� ��A{�+Ʊ-�b-�pgd�e᳙}1���k�_�m�����P̓%���X�FX{���z �$,s���L��u,��q���w�39��Hz�P�>6�*(l�-��4��R�^�Td��JD�]�R @O)H.jKw/�Sk[}J�~�acp�A�t��V:z	���є�%e,� �ۤY�S{���6�M|a$�/�e��y��)�W�&��R��&�*
㼝�Lcc��:L#��Ӥs�J��@�d���p�
�.�.��H�g�|�!4?�I���?�Y�4��?|t�����3�^M"�B[��\،�4�^��8 2(>�rg�G?R�L��Ne��Yr�Go���N-�T���Ӵro��g�O����"�,�W�)C*&�u���K1�9g
;�:����}�g��d�#n�) t�Q��p��B��7�����99Z��17<���ﾍ,,��D��˰���vZ7(�W�;I�m
�w�k^�4i���+�A/u]$����ȼ�C�A�W��z����y�[�[�I��VgQm��M�Ԉ`�l�4����5�#H�܂e���`fT x�T��'�[9���7	�BO�bq�9��1��´o����f�$c�/�pۧ\��1��K���d�l?�kf�i]�����8H]�.g��#(�`�d��&q��K�^e�T��_�_X}�dcm(6���\�Ս�v~R�S��t1�/�B��"���ȣ<�Ջ�&��P��a��R#�q����`B��rQ1��b;Yd\D�O/�)`U2�a��e��G�e����I�$�>P;�@��,��ieK�&�?�BG��$�{`���߾q
�:��T9b*��mx��=5 �/�������ŕ��	��)+�p'�9a Xr����7��65%�ȈHx�K��h�<Qg%�TS�h�F\�=	k�>Ɏ|��'�[A��������b[h�i ���B_�/
X��.c�sT�-V���rM��U�"`ө.QΤ��A�-���23���<��h�Z�%\�"��Y<ߧ���P�g;�"�/f���0-t�3�p�e]xn���0� /�=�;���N2�Es�Vn���rj��qr"�]2���1;o���Bp�X��wr$(T[�W-GY}o�VS i�(�uǤ��}���h����R0��6q	)�-oVK�\�� _���9\�@��b����S$��AvoU� S��[1��������#���[�=�� r�m���(�Nf����I�צQF:u^!�JI�\�iv<~$0���k%s	��1ٮ8��aݹy��ፕo&1G�f:>>i�G%
��u0�D��1F��Q���<+�'ŗ�pl��&�L1��C4�.N�)9Qe�|�����dʹ0Am��6�[N6��AޘJ~���^Hxgi���m���Կ��b�܈�	������^�I�R�t	1MX���Ԁ�9��pn]���AF�����	~�]�ķ��o�Nx<��DrG���L�:���W����G�w+d�*�_Wo����5t�d[ݯ��ل��螝\n���>�IC�f��GF���
;���K�S�I�U�� �*x���������&a/�t�7w'A���0�D�^� �9�[5���q��BX�}��ݛ2� �*Nx���i��F�p<�h�/��p��Q4�b���w�'��H2����^.�[���͒�:5C{��L�t���@�H�ǖJV��O�S�˺T�~=�г�EuQV���^��ߦ�ȪZ�T�a�3)i���B�\*�}��j֪W�/�̚ �7#ոU�c��VRS��׼�uY���a��$U�@R`?�5�m�����KhBzH,U�v�fR}�5�{$��5����db������������za�Y�]q&W��(�i�"/�]K�A�nX"�s�����64�HE�ݑ%R�!���x?�K_��2P���+�W���Q�������� ,�³t�fO�Vq��$�Yw�A\�"S�e.d)@.` Dl�.�i�t��b�8��.uB*)���tǛ�7 ��k˾��)�y�mF �:Zr�h��.�3c�ӏ�qڔe�B{��p��lhL�_�k���q֌����R�0����P{w�^�1x��؍�?z�)E����h�w�[0��*��w��0�KlIs��Q�B��5n��
!N)U��Tb��*a|�/�˖�� ��%��-KuUY�����u�H���D�q�FCE ?<���R�Q��J)�_���M=�l�TD�t�ʋ�!�������P4-�q6���t����ǀ�H?�����va��[�����L���gF8�ޭ)��#�Zw�Y��y�4:ߘ���٤J��=g�ь$[���j#�BoF�N���	g�^��/�r�Xt�hD�Y��#����}2����c<�+�;;�:e�c�I^��HUwyCJ��ʝ�6Zx�Q/���Jy��f�� 1�$�L�H��5�S�}�q,�-��"d���m��w��x)^�9�ꑓ�{���mĸh���Ln��
~���5��oE��t����xCܣ1^�����U*��HDc4�j9���ip;�޳)G��8����)���V�R08-<���ϡ#Un2.̾>5��¹�v�I�I��w0�`����9�i������WRD�D�����Ƈ��F�I7��P%��o����1e��'zԽ'�}~�B��3�ܴD2zM+n���rm��dI�r��|A$�T��a�i8dv�e{�R075��gL��ɫ�Hv�y�l7���"���/��Bo���&�R�)����r^F��oҷZ`v��s�����<�>�����x{�����"d��{C�w�*h���L	m\�	sm�h�+J�}�K�����]"��nN�P,����J6YR=q۸�R�;���[Uێ��A�h|���дll\
�7�g�pw�bt=T5�rG5->�U~�'
oi��	.Njt�>r�v��'��4�V�H C0h\���`4:��'(��Z�V�#��ɋ��i8$�2a�PC�G��P�0��c�
���:�=ڳH��Q/=����1*@��9
la�wS��9�ۣ�tˁ�H�bc~u*"���eD^4�LoZ��3�J����1��0ph�2���gF
���ЍX4���4�~����R3x�ۗSd����Ne�z&f^����ˋ�0	f�z���c�/�YA�BG�TC�%O�:)H��|�7���U&�cG��R�V �}�]^[��ԇ��8�������w��ҒHD����/��jo��	����x��3|���ɻظ��Ϡ�Q�u ��Ѕ�ı���\�^�/��@��p��m���#zj������g��`S����:�Ѯ!Ed��h�Cn�P�F�������Y�T3� �����VAAUL/@��>�rr�/�&�[��n��u`�u=����@���.��\"Щ��:�5�T�9��B`����P�Y�U��Fc��ujB�\�'
Ϋd��T.ӈ�4,U��l��i���Za-m#;%Q2��<MQ��wX��I����vlN����q~���Wm�t�lI����|G빋�u�Ro�� ���̞��R�O*/l4�ɠ�����Ns����(V�8���H6�l=����FP+6G��ZG�A y���U|'s��$�^�ĕ>Q�h���Q$�Kz).V�罁��C��qxW�nJ�AH�Sm�:0�0k�ܵ���iTN9�A��m����j��=Gư��JR.���/Ap��|ů����`h�C�7��&��S��x"0�|>�Ą��uϱ9 4�{����PVn��2���Ma��#�L�_��^�!S�D{���+,N�v�nImm ��5�{�u6m-
�"��|��B��õ\,���X��x曎�DB�	~2,�r��d4�������nڞ��umcn-�(�R5yw$�`�?2�Z���v��@Vp��,y�w�����T��Y��krl�q�J�H3�@�|��1m��B��<�X�T4=W��'¹��Iw�`�QY3L��1OF�������}��:����Z���󥖩������󘛐��+��"t��9�3@�Q`��S�zo�a?�')���R��ҮH_�K�=SW\`�>�  ���y �O�mlTA���pݥRF_�?H�'�U{$;�4��W �������vґ_y�=����T�� r�ɉ�:���!m�RxJ��#���4��D�t����LL�/���\ �-�-B�����p.���ۚw?��9�=m3���fzRW�������>�N�-z��)��:՚ףK>=w'����}��ޗ�^�?7���q�YB��'��ݽ��HZ�\�� g�H#SMyn�&@V�?s���L[��Xa����ޡI�>$fQ�e���t��G���F���>��N?��3�E����K[w�Yx3���D���������&#�1ő|�#@����&14���ed&�=奡sM7��m)O-���{�6�(�N�h��Ld�cPN�3sScp����;A�� g��IO ����0n��Q����_���H�u��=$js%��.��������jF�\ǈ-�z�ʚ�s!�(������:=�W��z��c�t~Hf���j,��:��&��>���D���Pu]~ѱ6N�K*귂k�v�^�0wi���JG��*����nxz=;zѧ�@�=��@�E/0��I&��OוiRC��CN���F��@��()��Aܡ��cg���Sɞ%�>�����������;����k/"-#]o���n���v�`{E+Ǫ�j�d1�Z��Ƿx�����>��˘�oD��?ޡ1'#"����K%��^'��N6� 7�������y鱣2�:���F�Uu��k��L�3Q0`q$�]�K��&Bv�k`wsZ1ݻ�0��e\�m��0kP�����$X7�u1:3om[s4Q��2�&䭋��rO���%t����"�~���TD�@�窛�]�F
���F��w߳g�fFXH�`��cR��S�C�)��4�N��6�'�<�73e�qG�W+������%?��D��f�fE�0��T]��ؚ�8bU0��uHf6P���x��j�	�<�k�$�2 �t���H���(q��\�W�1��ن0�j���2Qe�n�?]�(xf#&���auR�U���|g�_����:�r`̘<�JU~�iJ(>�)d��
�E8��'݅�2�O�K����8���"W��a3_X+����%tn��m��+Mf�D%��$�O�o�\CSp��&
��v�W�"��/����,�$0Sjr�/�����������ٶ�/|V��ة��Т�������b~�g"��� �A�H��#�:�/z��LU����� T0����ty�/�Y���EU�Ǳ䣖����剙a��b�����\���馺͏�W�εy0�]��7Q�j=��A�cw������ ���Ƅ�Y���,�S�)1h����^[�؄�F$��TMV�i�@�,�J:�P�3e��Hv'��
�;� �&����R6�����1R5D@g�D�t�d���ñq�P�;+wp�^`�������{�*}��M��U3�bm��ks���;�ޓ>�Z<%-Ǝ��$�����>Q�;��	k����*�A��[@j,��]i���� �G�al$I�����M�]�կè��cB��x�;��-���@�m�rU����X�"Zݜ�����w�H�sMF�^K,Q�p�D�&L^��������W*
��wR��0|����u��`Oq|a�v��#%��e�{�꺀8�a6��%���xƏU�o�惠��/V�!7�~�I,�΍ޕ䘻���C��c߳LA����42�5"n"�"���?-D V{��潦��@ݲ�d�iN�U���(�P��<�6Bg�ȡ�!��{�P��i5^��Ŭ�X���®#��h�\�/d�߉>��FG�U��tB]-����̪����M��PEAh9�ITځp˞-ҧ��PDV�� ��F��6��߀���A�4���y鎈�=l�`6@
��A��%$���j�G�5��6N(y�����ڞU=&����P��H$7�����[�Q�;Њ�$i���L�ޒ݈�-kI<��!2m��<�0�b\	a���(<u�s{�gYI(ϑ��NK�,j�҃e��H�C����V�R����@D�|�
�f���I�B�'`�Um��#��,�oָ�q����vK��Z���(�2Ty�ca~�3��3��Zȥ8�#�8&$�
ik��ޮH��a��gK�\b ����'�S��]�f����$G��V��:������~�w�{���0�`b��a�ZV]M�<o�L1�˧J��R��hR˛�y�u/")��
�օ���+_�K�7�/�I쎬M���{�
��lL���0�d������|���0)g{
�����,�-�
h7�;������1��9,�R�,vxn���ĥWa�bc,�}�uN /^�-�_R����(��f��Zr "�jH�[7��%�0��l�ozh�
��� ��.�G���
_�Cv�a���L8���ސKc��H�O !c F�J~#� #ch�`bq!��_�h�z}
iT��	+��ח��b[{SI?ϥ�*�E�����b�r�$�CH=�~��?[n�u|R���̔�a��5�,��H��)̧�Uj�7����N&�{s�)& �&6s��u`�}�K�:G70A�_8��ww����$�!�*-�{�����4DԨu��N��Y鉁��"%K� ^��bO��2&��̌j�<�:�Ku�6�n��Ԣ���|^�Ӈh4�Wi-)mw,ꁿ��Ue}�0��[A��P7܂,;���y%�?�P�~2��^R���u3������f�P	�c��.@Ah�8����m���oB�q�9u/���X2�(�s�P�Bۡ��0=�5�"��]����)P��&�,\��]��ILtE��ߦqe�q����! zi��r��"��K�F�v�?�Zʨ`'�'2��6ӳ��fbqnqV-WW_u�p	V떪����m�P Ŵ'͏��n}C���d����I���Z�`���J��A�~�N9�f�޽A���ϊ0\_���әo�s$�Wy��Q���7^L�P� ��[bf��\�BR�l�����6�B�|�:tV1�MG%znB��P�쎛��-pO�p�[K��~�E�=������%���w^�2�{�;8t�^nxΙ��"��^�����q3��ϴ�M����/d�y4A�/�ʚ0BǕ<��G��9��!XQc
�3�$�oi�M����p[;pR=�m�'�{=˸�!t\h�QJ$�l#�����������@��2�u4+�Fߢ򘂦��YN
I�����+t��u�Oo���n��`L3��Wn�}X���%��3�v5@5!��st����7��m�Qj��5
�=ʦ<Nlɛy13n�p�`�NKJ�B�A���j=N�5F��V��GN���2@�N��~�{��L�=�V��K� �C5i��2؃"4��PL���q�E��*rE��)F��E�W��kݓ#�����c���S��y��
d��3�ŃZ+wŴ'���b�Y�-�7|��&V\��S&ӧ�յ�sMP�'h�� �`D��cBҒ��u=�-��n�(Q�p�G����j1�l�፱��qd,]{dH�: ^�{�l�ljL�NS}�|����%�媀z�y�D�$*O�����_}�R�'����}�ה_W�Z"�T"`~���4��|��S����{�G�A�-q4��u�cDA����;c�+y͉���P�&�7���}��������i�ށ�hU�|����Ͳ�h�y3��m�M	�4�F���̽5,f]7M�A��Ĳ�|da1�q��,*�%XC #��'��c:��?�QG�H���z��qab��-��N���.ؒ���I�e���n���x�N�i8Wת�W����N6<�P+������_����wj�S��h%�b������5�Eq3w�& M{E�����y�J:�-��n���R�>:� ��D0 �}H5��wȸ'�{���>�Nv��J|��%��z�[��#�O^e����,����d�0i�,�o~d��Pܡ��J��C�p?;��{S�g�{�j!r�Yr��d6����W�5���֋���4-<y=,؞��e~[��\ֲ5�5W�]���H)ǂ�%���#�N:�-��4v��87<3��ғ:mx�U{�9���$�Ǿ>"���.���1x|F�l��L�y��_'����>ug �m�+��WO���p�����H<02W��o����rć�#Jt��rd*��D��&�䖓�^�N~�B��U������8�*x�y�S�Zq�3,��+���Q&�/ՖNr���^`(pۀ��<(�<�И�_dGL���k��[�/���`�^D�`.���[S]s�-xb��tNB�>"��LyQxD��v%��b�����y��d��N�Zx��ܯ@R'�����a��#���c��ҹ���ZbEyM\�o�B�'���oٛN/�l�3�?��;�t�PK[��� �^�#d���D�L	3�ڟZ��w7~d����[�v�<pʣ��#���B����#�Ҵ&��)�)$����IIB�oiA{��e�LNo��x�]�%��!��~U�,�
�kͱs�|o\/�<��]	�M^���ݛ�ʗ�����8�0�� ���jOǶlǇ$s��E�[��m��/J��a�'*����~V�DM�����`c��«ҘBp	�	��E5���mf�F�-����k�yvy%^ai0�����cd��ym_����R����޽UpmD%��F�c��xCN����c�1 ���E���2���\�h����b���\N,J�᲏����l)e���ʨ>�0a5�K�����>�t�u5����,���A��̺OTs���q(�zH�r�B�ÿJ� v>���d���b��]\��^�xNs�/mW�_�DZ$+\�Bb���_�a��(�M�@��U<n��n?m���6 i���p0z��äXNY�����8�ײz?�D�[H�e⪻��JA�&sO:�A�.����ͦ@��7���E ͖ٻ�ꁀ��t~���
?����}Q<[��h����P��f�S#}C�@�g!$����sx�a���*�.���us��!��A�]�K+�"i�!��O�N,���X.w�\޽r�i���Tn�Z ?�[�c��uO;��ּwUڌ�YO�RVG^O�'F	�}��M������}C`�:�=��ʞj�p.�N��퐦O�DV�����#��ѽ�Ry���G�)L�Lb�şsQ�H�;,�y�S��N�����F��>�g�e��mN���R}$gL��d�� �C<}�?	$��d��Ü?O[:W���Y��B���߫�T��)��6aP�s���ur���t�7FP�E_>d���W�v&Da��𭫎�U�ڋ����ع|%*�����޽g�x�hQB�AO���[�I�-I�@��1���՜�5F��?\T�t�hRn���r9~�[۩ ��E$�����,����ݷO���@J��R�W�T��M�hʊſM9�9�
�����BJˤJ%7Y�~�'9X��	Bz�OT)B��=�H��2�=�Ο0�������iz{ocr:6�'���=<fIC��z�N�0��X�F�P�w#�X�5Q�-���)�D/�#���/�	���ϩ�7*v��z��m$N���bŶ�^^�L�O���5O�M9����@Zj�J�6�{�%s&�2���5�ى���N��Rڤ�s�r�
��5�Ǩ��XlMɳ���:��*��A�Ɏ�td��,մ%�$=F$�����iR�&�1+ܿۋFU+����s�y��7={�\C�|�%��3��n?B��3ݶ�[�eP�z
K�iFAh2�G�¯*�=4L!����N0�>�(�x��(����!B�=�`H��`�_���T���b���-����m�!Fcv�P/��?ٯ�.Ã�]�@�u�Y�O�̫����;F�Z\�b�G�+lRE�&t��5y�K�,f6af휅�ס*�Q���K'��������Ϙ���Ղ�5mr[��׭��yPP�Q.H��Q�������j��K�8��g/��=u��Ǜ���@�G�w�O+�[o�̈�x
��3�?܆��{Y:HX'"�:�����
��r�`��`�XQ��K1�W�Y�6ÂȔ�ޙ��e+O���W�M6.�l�к�¸����Н�S��ؿ-�Rh/ןQ�1y@�#3�5Ŵ�'<]�(踂sK)A�FZh�
�>wKPeq*�(�'�HC�d?�OMk��a�	Be�!�=�3��ڨu:-�s��<��t=�5�CZ�vBKi�Yե�9�J}��:U�`'����E�nqx尞.Nc"�BR��r�y��kx�~F���Zi�V�Q�$���o����ܨ�2p�5?��<�����V�I���|֊�2
v��y�E�P����O �yo��S
�e^��@�E�%Q�C�fS`D���XWWq��h�٩��]�R8X�^�8q=я���A�X/RH���]>�lb�_A�W.����s������;N/ůdyQؾ�����'�o�ZdU�fc�K�����ѹ�,��������H��[�q@>�(t���|.ef���9)MxV�6�j�+��|���[��j���0ct9�a��D��G�R��iG�.�֗��W��_�b����zuQ ��^K�g�t��9*ň?{VK��X2V��m��(�LN�=^D+���u����H��>l�e>xI�B�#C��p2t��72u�*iq膌�Ԃ翡�4�b�p�,��*���Ii�ag3�-�G�q���O��P�o�/��)�E����y����y�	&�݅��rf�?t2��;JD�bd��7_^��1�CULC	~�dcW�K9dҹ�(q�?����aZ)G�M�ˏ-�R ]-6��L8�����9��0:ĔQ�:� s��/%��-y#�w6H���r��S���:�FC{P��< !~�r�{��7��8�&�_Υ����b���0��Scr����SAG�ϑ�J��А�@�( �l1̸�1a`PH�	�����/�O��dui��ǐ��	'y(b41�����9���#��3� G� �e��x����{mك�1����jT3(��X�.���>�I�lm��X8�i�c�P��Y}��dYf��C��B����b����8�"��~�É'�'S�/�hM�W&H2s�*��
3�,��7qM+�0�H�Ҍ�s���Ĩ�+<N�dg|Q_�0+��ӿ ���s�!�R �܀�tu5��H���p1�L)�@�a����*F��x,|vEx���ʴ#P��
Ezσ��UR�M�*�4�w]��-�G�UVև4�2� �:P��B)["��Z�BN�8�m�~�{��R��`�'�L����-��0,�u�\�h�ȹ]��4��i4}-t^�Eǃ��tt�bO@R2<���آ��əz^��i�
�k;�2�����:��Y>��Ye�u{�Ǐ��r���DE���dK���Nh+�+���m"q��{OT=�7馩�3��:=����ô�E�������z5�A"]Ȕ�{ �.������"
�k����+gS��VG��Bd��[�0�*w撎��Ǚ����#�볂��J��>"����?*�`<$���Le���Ѝ�Օv<@]4gY�捯��0+Q}+Lj�F
�ҽ	DB�+���4�e2�	���y{x&��9�:��P5��a��)%�was'$���ڡx�-�֞�8�%�Ej�'^ߵNeq�!\>\V%S�tw�Аε0� ���{`m�m�%$Z��OA�F·���~��\f���c#�U�L'݌�%ͨQ�Zh;{2�����L�S+�����r4�Yv+e"��G��zZ*yN�B��0�Iݱ��F	ב���}9AP�����|
(�v��ĸr�I�1�b0��(`XY�g �Z�u!l�T^3�PM���t��[����29B��c���,��K��
�d��N���gm����zT*�q>�W��߂��I	f��"���\�Ǹбۼ�V����-RR�a>�e�ھ���S����b�x6�"V�왻(��E��M��9�2�B�:�mx�.TFtN�g����a�}J��ϱ�z�νF$
bv�o�h�`��)�i�sXe�)�|p��3@&�����m�?6�i��	�D�����DE	V�y�'�n�*Qk����[e2� -gJ#����.��pR2�d��㟩K�i��-ƑŊ7�]-~8�{����T������@�Tr���$-ӕӶ@���=W����z���ӓ�d��^\9�꥟O=~��:��7(�7y�Ŗ	��V��`1?��S�/9H�I�lDv}�Y�����`�є_T�m�����i=Oт`3�ޱj{��%�>�/tA	���I!�>�RCo�yW;��
eT⢅b�����߉o�rU��2��
��5+.����~I�^�^8�y����~��<�rp�D�[8�X���0�;Ei��4\�/6�(���k�}Ö����x��lwA���K*P|Yl����0A��.����DN)�o'6�p�s$�I�oj���w���q����]�n���`4S&��	�I��ԕ��JX�
��G��	$3V�a8,�����c��KL����&n[�V;�2W��z��~�-s��ߜ��@*�`z�c�0��Xg���+ �슜��T�P�Q�Ho�ȭ�1R%�Z�u3K!����̼�U�n��+B�����T�Fks028W�}]t-H+����#����KiׂT�q�n���UE���f)Z,6  ��"���� ����ިOJ�9N-䧛��e���ꯎ�޽읜PA>��8Ds�CW�=��IIc��5x���ހiL��O&��
<_4�JBt�H�'��N�@N<��YG��"\'W`�_�H�߮N����9�#�oD��� "+� �_س��i�G�2)}��4�Lt�t#9��ȅ� ��?��3;�����ۈ�_�ǲR
��O�7�ʐ�h�N�
���O|)����Y��K�m��B�Zۻ�C#�E��r�E�[OF�'�ܠ
����p���h���+���`dLV_�<-��E��|�ٴO�5�������4�$��b�k@����C�H�~����J�[�)W�-��Bq����I��*�(��)����~����ޏ���_ ��%@�@���N���x*c)�-�$���6f+�2A�5/��A���sRieo�1m?s{P�2�Jv�e�@��~)_�Q��d���0��R∬�3���RȄ���!�FW ,L��si�ʊ<����v%�іx�ܶ.�{��E�>^���R�H{ϒM^�4u�_NѺc���]�D�T��J���#H�PRО)��^�H.B�ˁ�~o�[��c_>�&V��"�p���/x%��4�w�xz��U���2 �ŢwG�I�{�ZU���K�:���[�����=�H�W����8Tr����}���$!	��8K���Y.E�n�^`��mD�]��|"q���Kc<��úG���=��I['�P�<Y�j����c�#$��v:v`H2���/pu���� ��t�%�s�@Bx��{2�sM;u���L݌.�X���k�~Ν*�Lr=?��%A��*ۮ੓!=s?�J��or^���A�w\��\��i���L����f 1����
�c]XO�3K�`�l��~V(d-j�_r�V����:H�sB����[G�F��m d�*#��
7�ii�d�P��^��c�+���U[q{N'NH�� �U��;��mP�l,����b=K}�a2qM�
�e���,���Xxo��4l���=�����n����~��K(ފ\,����߃�e�ѹ��r��
�㩧� V��/�ݠ�4��{L�m�w��LG�c���*>k�v�?��+"�x�C�z;s��Q_�%[�`X�C#�a��
�w� �H \eeE�f��4�\��W.�.��)���j��-&��_����՗�+��RC�_�4i��w����M&x"<MW��)��u���M6Q����X�}�Ӆq�dlp60�)u�ui�
P5��Q)�����s�!nK����_Ѷ��lz�ǣ&'z�g�%����ś3N�4\�8űS�t�1��]�V��#&D�'�`P���w��S��3mc@�v�+[;̹jp���`�	�
t%=Uy�f�ܛ�%R�p�?C�a�d�+�w��h�$�#�Lۧ̊7:w��@s��A<!P�pɭ��Ւ��2���ȓb�-����v�A��O����U�� 3�0lʃHBFBqu�Y>'F�e����J	���_��^	�{"®����8������i��/��&~�?y�]�7���nGX%�Y�
	n�z�w����窝�.����܍���eJJ����Ĺ!q_��S����_Ylkj(k����ٗ�x1�5����!H��!�g�o���+*VctFa�w��c�l��;M�cC<�QH��Y�:�L8(�%Q	��z:L�uUc�!�W���[/G D&�8��)4h��v���f4�f��)�P�,t=�E����X|)����-��Fu�6��\�#�O,��5�,ڍ�,q�
��ƣ�-��03 ��#�ʖVMg�o�2�f�8k���6�*LN	����w�C�;��_	���Y�ƭ�?(Y�\����2�}��}�^��M�?��h����Ώ��8�oǮ$��I�����	�4��5���Al�ݗT[��t�+�� �<��Tj$Л��vn�����A��7��6�9J��OZ�a��R�g+�[�����#�t�<<p�ԭT��u��f��WF�Y����7��o�*"O�V]���E�nn@+��j��Es���zfy�o�_W�Yf$������Ŀ뭗��#�8/���>�nG����t?bN,@đ��'��&b���K�u�����r"UԽE~�(����*�S�5C�`�ȏuTz̾�0��<�Tf�Ga���=�� P�MF��?o���P9�HX�B)>ꢒ��=�줋z��,��
v���h�T��X˵	/Ї�\������/.��wƜ�2��۪K���E� ��vRx�:�F���"By�F.y�pj����"r28��@�`̚��f�d{�2��xt����	��S2Ǜ���¼��B�����s���� I�#Oo�
����P�K]����)��e�_N�V*�]yA�vݣ��k�ܩ��/6�tP�������M�*�f�R�bJ����{�U)]nW�	��'��&@�r�s���~�m;�i�,"�%�*&^>5( #�v��.	B�1�'��a��.���=�b���{Uj��%�L�Ƌ����Q����$�3I��+zL���	5Z\�ܐŚֺ�w뵍�V�r���B��q����[\�-q�։�^��H�/�_x1�[�:��,�~v|�a�F�KDTL�l �E���qQ'��1�Q�-�^hHy���`S���u�1���,�j�nu�b�� �("��>��ʩD�a��Ϻ(+����?�̴c�ZT�S ^ �\S��ut������ơ��j�[�x���6MI�:�h�4{{�<f��6�wY�
�~��]������H$P�*���zSq%��R�OV7VN�bn4�	%�Ѕ/q͑"�1��A@� M��^d�k:��2N^ ��ڒk�`�.)�钬v�� #��}�E /C�zf�&�m�*�`�	� }��F�?���K����3���#pe��ӡWU��k���-
�VT���mj��ZmJ���p�v��6�Ɓ��&L���!�nh�Q!5HװD�Z���w{j����2ɞF�Nŭ�����S��������g�)}_9C���R�tY�]�S�i�o.-@-<̊� �j���zi�b�
�Aw�G7w��ϔY�>T�����x2#d
k�Ʒ� �)d�cɪ'&�=�9;��Q�v���:�t]��ݹs۶}�ژ��>_B��{*zM��ٙ�F]�s�1A�G�o�k
�0�g��:C�S!�qg��c�{'���tx)�\([�FR�C	`
���@!�D@-����ie��G /r-V���z2�t��A�����t`6T^�����u��ܧ:�&�[y��Bhb��6h��Ȝ��(�;]g��ë$�0ݤA��h��(�r��2�
ϩFD�6f�e�Y���=���L��ܓ�mD�����(?��N8�Qɠ�������̲��1[���e��VW�z����ka��Fx�k��|��ވl�z�\�M�\�_���꽥�*�Y��q����֭�� 4Jk��,�T@"��S�\D�Ы�}6X��٨&ket :�vl�e`F���1��?x���Ɖ1���&���>k�$��i���Ά����H�3%�{ �����{H�ù1�4����g1	%���1GB�H� �e?��;+5��Ǝg>A�Dr����迥i&��&�f3��ŀ��1��?zy/l�����^+����r�[���#���`ސ �-S�	���ڋYRݝ�j���j�H�����t�8�C����
C��,Eξ]��Q�.��I	�/���[����?��E��;CÖ�7���9V<�	o�Կ���VDFt_��3�rx���)a.��8{3_|yG��wCfjBS��	['�����O�2�����I��v��
3$y�ܼ���Уa��^Y�0� jo?A�٫f6�q��6׏
��.Z�cu33�2�l~E+�40O�L���,�g|�xq�֦Mj�c�w_|�#��'R��!?{�*�x��
�~p������ے��o����sɅK�b�a��eݒI���Vq�ꖬ+���	��ICw��$-����-�[���j�޽�n�q9����q��[`�����uj���`|������Wk�7Ҧ�any<o�|��X�2��:����`�5���^]�x����¤�}|�!L�_��UrLk�5��5�n~�2����_A$�{e=�n"2A�e�_��ZƯ��_����$��!̲��oo�"A��uF�%)�h"�K�ܯF�����3�T�J�ƚ�m [�0��h�=FnF�8gY:�r�p��n;�fK��P����d�Ñnļ���-~����.:	��eW]/��vݏ�]D~�u�2Y%y+9�)o���+ۦl�`�e�v��21O�ش���ɸ5��JA����D�}ˡ���v�ܐ�@6�"{k CEmcG��:)� �Re��q3�S
<ޤU��(9�j :$�}���m&B��:�5�7t�_Ϙ�d�m���}E�����Tv6�Р[��֌�{����lS)�ɴ	qcu����E�@�=0N���u��[$\.f�.Y��bA~�>�47�n䍘�����GK��A�>�Q�����͖�}�@�p'̶���d5L��AK����G);�����<-�x]4(:A>@"�G�g~K�$'��0���t��ɇ�m���G��`.�����S ڿQMj��ߦO��I�U�$�ѡ-{FE�Y@M�WX|�1��F��쐑H,δ��f��iB�R��)�_���=⚯u�+�J�~����w�>�!�C�+A��p>Y���ky�#c��S�--�� ql���W��6��Z��������i� ��C=�v�_l"�8���̒p��/�- {U����Z,��/Vݕ4@�PqF}%o�bgx��M_�O�ӣ�bq."#���=�tI�����D�S�O�DA��{���X�| b���V)i%�8�Ň���NP2I/���4�>�h|\�*A/���P
T	r����D��Z�!H{�_�EŠ���̷������D��+���m�=��)kA}4|�8_`��ьj.�F7Ӂ��c,dJP��ƔH�}4i�Y*Ut�I=�j���\�ILq~��-��²����9)����y�"s]˼�n��1�W>��:��%4�"Ǖ!�L�cH� �Ly/P�Ä��7�5O<��H|�i���GrSW��\I�������dcf�f%���m�ۑ��ۤ��b�<��ɭPM��IErq@��/��ہl�K��������o�Z����9y�H+�n�4~@Q��X~|�\čhN'W�4-��	��<Z�R.��%����^�g<��Q��_n��P0���g%�fC��ҥf��\=/8����7�_��@IDSI�B��xz������%��^PEH�z�=x$�f2#����u�C\�_�L��·����T��H�+m�Q�	�n��%G�-���������	H�mSÉ�R��{"	�\th�f^��f;��T�c�]�sf�Ó~\�V[E�p�4��Ѳ"j<�\�����#}�[�_���(�N�AJ�릇Ҍ"]���o>HP&G���n��� ����x��)�]r�_���,uΉ�]��񜣨� �i��l�9� ���th� �Su^uOkM��cAD��B������h@���ɦ(���F����%HAz���A��1�1�TcL=�r�ƀ�_�u�D�klDN����=�M�[o�kV�g�87f@�6*�[�¢�T3�^���� p !F��n�8B����	o�q�swț[ 8��������7�p��d�	Lz�#�]̷�v@>�,�W�3",���|1����Y��lsϹn�m �U����,���G�Tfv�^��@v�w<>�o,[�თ���>.;zV����ysz�� M)�����t����g=[R��Q ��5���� 5
j)d�n_�$͙��	]�g�"n\�0�i��:B��0�re��w��س�������ׁζ�~�^�d�^عuvl�C���s�R��N͎���;8�]�B1!�	��d��������W䋑��[�D]�&��Ὧ6T���3!��o*'�q=�o��*�?l^�)ġ���E_'n�� b�
we���9e�]�����)9acwG�*�A��C̄���Xɱ9.[��0͇�N��A���C��C�mj@e�ƦܢO��0�����d��
E��L&�/['&"�Z��}��]���Ur���%��aE��`��#���P����n�5�?����^;~�,������)k�ABsg�]w�{�����u2����H`$��c:J��o)��-a)@�KD�Y}�7A�:�i��cUa�M�l��)xS�K��x��B`y��l��2T1�
/���z�t ����ӄ�P��~G�����f�]�:%��Xe�������+8��l$T��=3������p�,��2ͥ��Sz����ɥ ]�)�I���M֙�sY}O=�wp��	��*�:�uȖr��(l����)��ݱ{�X������Pӻ� ;^e�:N��&)2���TT`�19���}H�#Lyo<�%m20]�Ϡd%�"���K)�Bg�.��]��Z1Q�a�ݪ);5���Q��kW�=��P+�.Fh�l�f=kviI��J{���n
��P�B��S���ZP6@��(��k2��^�l�u�Ո�Q��g�PRV�S��;� ���,.��)W"����j�Y�w�F�w�>欒����<O/29�U��]���n��l7�6��W�-�_�G|�^����}D2�ny�C��9� �kX
5�ϲ��A�iq
y7��-��nсm��s�侚{��lQ4�����m5묪?�pA��Ŵ�����g��EZ��b^j�
�"k��� 0s�^ch�.�T]_�h��f�n��k�%㏤�c�#U���\U�Ȁ:�\T\�c߮��c�wq����`~g�X�
"v���VB�p�i+�{��(t���*��W]ҷ��Hs����� ƽPu��@j�|^X�鑈�׫&|��0�4n��x���H���+4yKQR�:v����I+؁�l6�rgT�es�ac$��$��*������.�u�-��۴?�����?p���J^�ɺ�j:���L�vA�?Ƈqk�< ��7�/M67^����c ����m�Ŗ��V�ٰ�����m�!��&f��MaiKv�k�î�Є�ب~:&��%u��f�1& QR����.�6�A̳7!��~��͊�IN�dh�xS�v����]�Z:��z�������\[�u#N��x��w7�o�������ኃ`c�E��>���l� �I��pJ�7o~Zc��ԛ�<|�D4���O��+����<5�&�=4Ͻ�����9[_��0d �K��9���ۀ"q+�ۧ_Q���'N���	�J��3�҃���0����Z�1	���x��4�y< ξ=�ܯ����Eɹ�c�I���b��whQ�9�͐�Вiq�O�CZ��e�)O�7},bU��_ LEؓ�v�<择�;�6���ٛ�?�|�C�yZ��<N�w������>�� �:߭��,���y"
 J<?Fo<�0���c��I�?����]M��J��G�d}�$n�3���ȱ�P0>�`�����c�P�*��PE��,E[a&!��J|ib�.�����g9����,R��v�Q�C<\���ᨺ/�3���=q��k��47�.B���b�\A���"�}4Y�6�w0Z�R\�Oh$�����ȍ&�Ou��|P��'r�ߛC��ئ�6.��Tg;nN��}y��i��pnF�ˣB���!�ع�;tԝ�6C�n0��0]���ʺ#`$���Y�R�u���K>c���539FH����Dβw��Qo�{��I��Ի	̹��ޥ 9�Q��TO�/P�\ũ�@,�@��Z�
��=Hb��b�{F�D����'���a��b�����!��F�Q��L�g\r���ǽ<�%u*�0��`�=ӱ�w��h��2��X|r%q-?�j5�넧��*�р�P�Dx1�Q�~I�
�%�R�%����w�\O&3�F �-u�7x#���Uk)�DV�&�_\v�6����2)c�`�����zj��o�j���q
�<�����'���F���+)6�:����_�K��b�B��tuܙ�i��*�Ϥb`�ѝ+��_�<�4�#an{ 9��&G��H�~1���H"Z��N9�E�E���_�.�P,�K�(�d��ޏ�X}�F���c�5D,����GG�W{�sO�����h�5�'�'2�gkne�jw��6��A{rm��:zC��J=v˫���T Х3;��'Z��GU~�5�M�W�l'��	�v�9.?��ز2���������_k�]R�@�,��
l!����qX94�|%}$���]4�^EKtV�!�š�>#vO�����x:o=��C.H�eІ���< C�5:�����ܤr!�?F[��b���i���f��S�7�P<�&.,�tɁ6��ٌ�fmf���޼d���YAߣ��QR�ç�0DF%+f�)�q��8��Nٹ٥�� z�/�Xw\�+kS��lν��f���p4�[RM4]���zwNְ�`Z�l��K�������'� ��!r��/C��R�-�����ᗞ���J��F�\K�+d����C�z;OG�sH��DdM|<�5��Q�	��,7jժ�6,�F�g��ג���1����#�6+��f��E��O#n�n�{Ʌ�Y�M�+��b�ڨ�vıu7Ԇ���_]7���>TW�����	#�j���+�?}y5"\���OZ��2?���q������傆��g� / �.||���y�xH��5n(Z��Z�;�2_v�o���S�>�G�Ysa��S&x��U��L�
�B�A�Ƈ�'`o�}�z�M�5���CF�iÚ[F�mr�R�)c@=҈�l?��A򫨘���0�,<������ ��C���a��'k���/���;w"0s����	[���:��Gt��T�G�ݶRX�B?����~kG1�P!)Λڣ��bB^�d�KX�k�Gd���LT�9�ㅦ��n1�T���ﰷU��+�M��_oS����q�·���rU���%����(H�����@�*���	/92�#E�e��U !�r�� �k%5�i���&}061�v��24�� ��7�O}��N;�'�B�/��� '����{�~�c�A�P2g�	TG�R���r�XEML�#5T$U?*�� �ðg�o�,M���]�-��f�o	I�"K����c�1:����0=��b�K̏�hok10I��/�q̄����WFR���EȘ\"f��N&��=[��k�^�p�h�	�u��B~�=�/�����{Nhh�k�y�Y��^#�O���2�	8�Br�\���
�ؾ�� ��w����ާ�ҥ2#�<�ݾ�@,h2l�O��]|d����u��S�YRa9�놛T���t��K*�r�4���]J_���3{�W^�z�n��7�|(:�r���7-�ܧQ9�$��xɛ����40�K'�Jۼc���5����i�oh�+�0��Bz���+�����(~��%��a�鈼�D2g�V>��- �].�?����2GòY���e�L�)8�)[C�[bs����1ɰ`�f�uQ�0vo˃�{�y�
������\jQK��f6�������M
,��y:}	҈�F��F�l��E)�ة�B
O��B4�E�Y����=�����I&k�'��D]^_hE�b#D�A�W˿;�r*sƸ�"r�����.l~���*3�����!/����ظ{C���^d�<�,�,�Dƍ�V�ɓ|��;��·eڕ�A�3�N�&�ق�ْѦ�١~{�K"@K�_��h.Þp�$Sy��������_��=1��I��I�#6!w~��Dh�$��ňzQ���|UL7�L�l\{�@݂&D"_�V�>�q��~��XTM��a�L�(����W���`r�����Z���R�O��U� wdI<2�
�%�ߙ�	k:����@���5W��=� T����h~1�N)+��G��b�u���9���Z`���Ru�5֐'տ	�t����z
�۰U��"��{I�z�O��>��-!��G�M�%��ݰ�u�	R�f���F
����=_�I��g��N�;	��u�k^��X�g�x0�ԡ+�AIyu�BHau
�.xq���z�>h��d��{j�r-�ּ���������{S5}�v���hMM�|CjZ~�Κi�����).�"n��o�����zb�B=�Q �9]_�$S����e�C;�&�LYS@̏E�ޢ����tVq�(d�]�1U�»'/\�ئ@m��ߺ��-��E��U8|����˓W��v=1��ox�-I_'
�,���� }ۧhg�Qǀ�;*����RDd���<���Rz�I-[WFD0���������#N��	�HX�8�=H��N�]TB4`�Yk�B/7�i���[x��2h�~Ց�g�lt⦙��0���,ný����R׌�u���	~�Ph?S���M<��"���׵Ϥ�d�R�t���\�	�h]^_8T���o8�<�&��$�׷%��� �G��z��<����
 �++c�ю�h�m��$����'��lƊ=6�[����X��W��ʰ�gqe�F�Ts��;b:p�ٌ(l����!�	h�t��$roӷ2	*C��(�nLp�u1� �c}��E��m>�2m&�'�+q�m� ���t��7�z��g�TvX5�HvV������S�e\(a�ȏ@pr�v�d�xҬ���}2G�2��f1� L���j�����F�q�R���Ft����Wg} �i+�B ��W���l�+6�=l��F3jt!9>�����.+�/)��g۞#?P���V��kL����߳��6aWD�����**<�6Z����H������ަ���+.��|���=����h���V����g0�*r#I���ݱ:ײ�o��`4[S ZЦ��RƬx�a;@���6��ܓ�5��nUG�K}u��7^�D� �G�d>��jSc�r�i�N��u�kuPӮ�&ՙh�7�(�Z��ޫ��	W��l�ɞ����m��l��6����JL�ds�V�t����"�P.c��7gE�y�V�]J����GT!�2<V6<�ڜ�\��j��e�Q$�/y3~�wF��fI�s��$R0���*'�]��f5Pכ�dZQ��zL�K�
��Zy{�DG�e(sTƮ�:n��SU�
u�%��0�O̞	5S����g�
�)ó[�p�f�g�+a�װ1�ڼc�@�6���y��*�g��|����$��x��?�UY"6(؇�)�
�M��̩���c �����9�k���Ԡy����gy�
ě�&�p��n��o\�aJ0�h��c�ݍ}�E��ۇ���W'��Q��7
��ԹOu_�bcǺV3�R:uFK���Vh�[5d7�_�=E�]dv�����!998�c�5�O��XcP�@+VY=���̉"��A�h�=d$���C�>V���Hi")HY
�٧�&��yk-pGF�aR���B��`���v��s!��24���"�/.(q�U�F�X)�T�m��(�����fb��j�S�
����N ��+�lnoZ�>/D�gyw}ʁ���������x,�MmX�%c�Il���s��7�X�"0�C���XG�~��)�C��F8yi�����q�%�m=Է��A����G̾�h�$����h2v����p��D<������}1V��_5nJ�$�L�\(.5KS�v|�fY8�<m]�FO�}˰b�Y����Y�݃t���ʡ��E �o_h��b�ӯqi�4螪7��9�_]��-��y(g��(�f�g�o�Q%� &�wv�)�˪������## �V/�>��Rl�B��]� 2
?���$%�/c��Z">�=���N���e�a����G��yL� ���-�NBP{J���j`H������,��#��L�uK��-A���5d����m{d+���׋�*��B�� #��������6iٯ�&� :���@���z��P7-l=M�_U#�e�����Kw�NEe�Ϊ���'�~�x�#	AyF8��;�P*T�
�%���K��[I�v��e�+֜�Fk�( 1v�;�$� �೏@�*-M����{�����K������8�@�.vg����"��W�@���6�}֝cٷ�w��1R��g̵چ���|?X<twj�9%��n�W
�{�C�=��-"�=Y�"��k�D��1���V�_�������j��U�=�	�ya��������+��6��K�a��`�C1���:p\���u4e�-�z�	�`i�|'�`Cx��D�3���H��n�xL�T����h�C�ͽ�	~��e%s��ϣ��t',Q�M���P�B�$WUZ��s�y�B#�rt�ϲ��p�1���a�Gk˱Oз�n�OF���e{5s 1��+n�$6|���(�EM���Iz){�~t���f�v�\P���!'���k.L�@k�i&�����vڒ���L��]��E�4���P��]�⏓J/ZmFh^ds*��f��ڦ@���&W���|�3�s~���+6p#�rRУ�m��_xf�+m�<р-zG�-��5���*�/ykբ2��Ry;����������x�����E��^�0C�k܆w]||�H@�����zp!w#̯CW��ߥ�c���bh��H�ۧD� XP�����������⥹�����{N,x�F)]��،�9�7�b{e"@�*��pH3�HtM�:�zg����e�Ƥ��Q�jb� ��A�8J}S��|- �O;���$Zu���T��'���pgQQ�"v��O�[]����"ֱ_����֗⥁r���O2�*N�L���8H�/r�ds!�'���}�Y��	ٵf��c,#�Ej���(�H������<9�2=&@�,+x����?��$#��qΨ/CW��9�o�"YPk��o��ě͑TUs�sױ0o�^&73���G�sޔs�^-j�����|��s�Z8c��`��ʝ�9�?�N}D4���$�P�W�K�M)n�/�=S�����J�4z�v�+� �u�e�]5�Atl��e8����Z�;�rz�m���{�_���a;��͹���� ���hwO�v�DB�ٴ�fE��.��Ɣl�a����[�+L��A,����n�1*�WQ1��3�B7�Ş���Tl�ǥ����`�D6��s�$��0�,=��v�Po���E�g� \[!�0��&�8�DѺ�LU/�z��X�����6}�/�CP�|�q+\��8�i9�e�� �S$��NЂ�A���H��G�cV��˴���_`��n=U_�6f����u�t�f%[��r,ߛ��`�~�`FJ6��H�D|[���r�����1�G�T��W�}�\���v�Z�Zq��1�n��G�� !+|�$"�m��i(�c��Je4�=��:�9$B����O(���36u�w�J�ҖRؑ,
�=��SG���cN[�4$Ʋ.���]Kv �,��*�%�xW�ԍ���: ����9Qi�,yzQq>
�|�Q��;(�v�Qw���$|�I� f���B�.�,H-t�8�46�D�&���"��O�G���T��9���{�o�?־e��}�\�;3e���1���θrZ�ۂ�>����p(t=F��r",�F��̭y8��a�M^>�h.q]���qZC_��s2�v�ݔd	���q�]�����e�?]����76w&d�y�L�'�-u�M'�Y}�[L3}bl|�	#��� �z����z������u��e���42���pAx,4�u������ʎ�"�L�E$�ۼ9�D>��Ř���L��[�}"�L�N��c���^
#�gi�]{k�d�61"���GU@G���c���q�q�Ħ����`op�o����b6��ɿ"M�`0%���]EW;y
Ϛ�ۿ���y6.}=V��Q]��;�ʜ"��#��˛����+��O���yR��+��{�قK�{���|�mz���O>f�{
Y������D�i���a�kK&8>`��:���?��yCź�E�QIQ�pf-���/z�F��gڗ�1�(���ߑ�Z��f9��#u�ESŨ�{��\�[��H���S]kP���-��byܚ��c/֡�#q���*���!�B�yC�I,�+��5�L���t�>�Y�	�l���k����ګ�q������ַd�ع���_qY=<FrO��n�������p�㲳�hE���Ͱa�w悶�(M6��c�%!��m㨴b�p�s��:�R�w��N0ǳ�/��3lE�ο���.O�������f��B���_s���!���R@n�,�;��/���TH�)�N�:hb�a,��StlV�G΅��c����.b%y��T��GN\�+Uާh���J�RVa{^�����z��K+��g5	���t�p�T�o\�eY:��o�Ai�i��	�����&,���6�^	�@ʮl.`�x�A�P]R�_���K"=[�9�3�-L Κӽ���� �����%�LY�O��"w.[G j���x�f><�qÞq���1�d��A�[ހ:��W0<�3��RL&�1�G�=���L��wjEgC�ճc��@�O�$�zqI��5�*��gD:�\�����s�nLW�m	fe�8<�4࿌�`BV�Y͜f/d "t��]�I}�!eqAmB[��B�e�Ĳ�̟9��L�c�ZX;k[om�x:J1@���4�s�e*��.f>���EA��}�k��Bx��w4�ZuDԾ�+�$��jtR�9D�������B��%�ň�O�-��pd\��i�n��F�Am�a�{�x-hU7z�)A5P��r���yW���$EE�1��7��;��E�=�����v	�ͱ^� Dq���y��HJ��W=�������?��Q@��n�s ܒc�SS�A�E��{��MFE�껅a���uշP��}�uTe�#��	<��5[%>�搸ekf+r�`v��W�!6Q*�$�:e}�`�R�a����r���u��9�O��)��b�"��wֵ=%�c0g�hy���:8H�{4�����w���#}=�7E/#u�Ǎ������"�yw�f=  ��Z�+ͷ�RV�rUq������j�*��O�LÍ^�u� ��M�`_
�e�d��p�y�]
S����n���+`�tՊY��y%�]+ǂc�"�p��N����9xʌ�'�ñ�=\�)��	!��z]��p�]�w��0��?uY�ȳ֕rkO�R׭N2�:���ؾ��^�)��)���=K�>��u⠯������ג�M �EX��k�W�j�5�j�����k�>��հ��rʘ5sIw��!��b��9��uLyC��A��)��E�R��OG�w.2�j��m*tyj��X+��!�e��A��w�b�E��.���H�o���P=����
=k�p�X/�hP7b9�t2rѝc��Ӵ�,
;x�	L8��
\�uI������jb�v=�nȦ���9L�v$d8�Yа��b?�RX�(������� ��ԕ(0NX�q��J^d͊�����$��B������}��$qk��Oh�JAP��Zӭ;�&FaQ��� ��.�1��If�������p���+L�+��뚅B��+�>+�1����\B����h���� ��`Ը���!W�LC��;����	�dP�i�U �f�9*:�%�&��Nx�yU�o�Fݍ��(��[�`���*��>	�q	�U0P�E1Ъ�Q�@���<�\�ߨG�Up����)��vt���਑ls�\,z�] �;�*�֣�B�d=�}�N�6RC	m;$����A�Q1 Z-�;g�,£�+^�͍T�gKIa�6�3;���z,���NF�n��kU����@�H�j6X���R����+_�-m�4X�7;+D�N풣�����;�4�%S��]�G}*q��1* �wm&�+�I�.��r�G�og��G-H���$�[�(4z���%ӹ��8�#�a����yï�z�-��	�Vq�IHM�+�^���}�uC�V@��d�F�Vԏ7�+�[��Off욾Þ�<%�9�!=%��\�/�����E�>g����WR���1,���/e\&��ё�ӳ:�nU�}?>�5�Y���F�\��d��,�=�^�C�;����s��pB
�寝y��+u�~� 5k���aZ�y���rgbr���:��s�Y�B=�	�}ち�jV���r~�����7}!}��u�� W����΄�mD�󶞓���_�Ǯ�[&�t��g��rP�>�v7w-���]�xc�~(��v��f�X|M�|N���4�4�*������ޠT�Ee������5��[� �[�{79�����ZqF��qND���R�O�ר���4R�`	�2�2�#Z='d������3S��JI"���v�YR�b�
2�JЂGy ����<��p6�`�	�s[y'=�	��u��&P�`y����p+P�g��h����ý��>�/s�g`��f��(Mσ�a�SS����b�����-� ����� ��6��E^rLd�X0�;Ԝn��'�"���j��`�%xw禧ME>	�-Z��9����1�g��]��9e�w�|�hQ�,)��#���9I�U�_�&�.��⏐KO���ͧ�{����c���l�E	�W�p�N�V0��?J���?�'�a�6ڑ�zնd!�	L�i�-r�7��Ƨ6H�&�;Sn����6�����vv'c�z���'d"�e�/S5���$�{��YLk�cw�3��ɗᗡ����(B���\U�%��d�A�b��w�=M�3ϡxGk���Q���,7g?t��|�?D�n4�������eT� ,8�j���Me����(ߚv&�q������e���lz���;��;��Gq�D��!ه5��܈��j?x�w<��\�o�/[)6B�n�2r�Rh⏖Z?꣪���/���õ��W-�rN*�{�ϔ"���1�\�r|�o���~�_Ԭ��,�h�%^:ਣ�ew��F{���_G���;
��38�2{W���ׂ�����$ ��	��V��Y���`Da���A��E�o=��g'u�H)�۶����X�ƒ��C���]e ���TN�h�;��2TD#�<IpF(��ݥ�u�A�	��TR��t^�{�����R�?`+��~��@��( 5�l��E0=�������:t��rU>��1~_�y��4lX��LR-���\g42 �1���3j73�rM�x�{w3D��2>Z<�;c�L�d� ;����p���5���t��G�.N�F�<����5��� )��p����w�ߨ���?SIۤ���� ���C�"�z%���n��-�r���%4���[�^t]e-�n4_䤒�oY��Ch|�����dB>�{.���"��;��Pv$��������]����la9��X�pAb����^$��d�����6��3���pa�IG�؁bz�5��[(ƕx�\�"�0d��*��6\j�sy;z��&�[M y�Xl\ �%R2r�;R}��s��H ��b�K��B7�G��6�W0��X�M�Rqʈ䒢��%Cw��e�����#7��vL���ն�U�E.LOk ���g�U��-t���,��ϵ����!�6#	3�'��]_��:�s�3�xQ�3��9l���=n�!�2���R3�u��x������T�� ����S+�=�a�r���<�9TĬ�
.�K# �6�~�"}���Mb���V�(b��!�*���e�"F���f��IM2�����ۥ��ɋ�!8��aGI��׹��(�b�FN��C��I�D��(K�+"\1ܭlH	�B��s6��W��@A]��΁�o�$�4�a�Ba�!ݢr<����k�f��^�q+��Ӳ�)�bT�l���Ɣ��Gt"���� �
�ʷ�mR�#Y�i}�i̤$��pi� ������s%�玶�h�� �p�8{�<�DP�����:o����L��S���p#��f O�'#�Y�Z��
A5�v�7x��4M�.n2�(:E�7 &*���uS�8����#�%՝�I�w4��+�䟘��>O�ƒ�%��.��0x_�{Vީ��x�*6Pފ�M��^��1�59�ArѮ�US�yU/�S0�H+u�c��������&����}��^��|чQMF�5˴���n�'��#vd%AK�1/�4x�.�>P�p'4j�;J��=PO�E��K�^��fAJ5�H��$��H\��_m1E���t{�<-�L���j� �{	ܻ�8Q����d$AZm�\��8s@5�*��Z��Z��Hլi���l�y5�r�t���3޽"C��'|���{�Sc0��w��^�իA�Z
a�����V�v(;���9}w�*ĭ�X�������>����;oy���6��%��s�DdtGhѭ�c�am��x8�tA���2��YM�4��hf����[��E�G������$���`��ǌ�y]��+��"r��1bx��ѝ�5)k�\J��U�}��/���V����gXX�4
�՛"��r�����{B�8�1��["���w�	��� ��VP���3����~O4��2-7g�a��W���Qrc�V�����U�U�#��m�>[Vp i;�ɩUS�8�'z߈��@Zh'i�ݵ��guC�L1ê!�W#7�T00�B@x��O�)I���Q@�Ţc��I9xlS�=FB�Vl��.�w��YSғ���W��yU9z���~�7�LL��#Vgl˷�ó֚~��Tҩ��x�H��΀[�4�V�wf�}���~��\��E9km�wI4��_Զv��H���0�m�q1Lr�Z|W�rn�-矖gIU�==WA�!5���ݔG��i�kVn{~nH�*��>��.������z��5���Z,�Z���~0\h'd�s�I�ԏ@RK���V`U*)?��J�r�s����v���tqcU|����I�؇㲡�e���rnh� l�Ob҂��je=��J���r��m�;?�R�r8�
(w~�-�X�0c� �B�IjR����;��`>�0*)]c�]1�/���_ظ��B_��l1�$p"�mD"�9�BYs�09TE��>�P�F{�E4j���qB-s�c���w���:)��O�L?`�Z�s?����dI��l�A�%v����2��#�R�X8˚���Y*���v����<��V�!��$���\q�r����Y�f����;k�e��� �(1{�YB]bY�t̺[r�*��m�����˗�9�S�"�
���tDo�!���%�����<c����jems�_��dX��ھx�w���]��3��qX�Q�fz���B�+�� �mz4h��~4�|TG�7���/6�s�Z��!f�<��9�m�l8V+m\� �x.aGCL�1f�Ċu���/���4�98�/s�������~�tI�\|�o:����\��؉�J]ݠ��#ׁ���X����p�;�[���A��#�1z/��[F\�9�/,�M�~�FLg�������frf� �%�͂$Nh�L��Eon��NC�̗�2�c6�P�nf!�Z�W��,���q� ^q<I�<V��z[k٨jt��L%au�p���:������E3�߱t�֋�V����k����zL�<m̲~X��{+)�y�&
���ҫpy7 ��N^Q:���Wq��R�y3r/ ���� |�b>N����ȵ��/�ym^;6H�iN�.e\j�}�|5v4�_��>%�_Ѩ�i�MJ�=BlclZ�_�.B�gCH��7�G����e�r`��[%;&��X��t�g)b��@�Mk�.��9��+K��p��W�������jLW�#!K�Pv����9i)���D��Pm=���9��ߚ�V�PW�P��0)&��~/Kǋ��1"�w�bo\�߉fZBf���`��-tϡ�]0�d`[ ~�T_�	vV��׬�q�U�%��S�e�p斮�6Y�7��i�{iU^"�D��@I�g��yn�Å����̅%��F��lСDLp��Ud�	||T��,���ѭv+ �O�PT��6��'1ə��3�2zQ�m�j������W_42<Y��u1PY7<F����,XI�F^��~����LM�N�v�8 2���l��JBg"d�� ^R�.���4u\��GY6��Y`K�@��n����}�_h�ĕx�c	���up:�L�� �<�Ĭ@
�7�
8e `\	[_jV����a�Q5c���4o#��j�Ү�����P�sT�1��w�5F�Y�����&���!i�����ø.���cm\ͅ�{����!����ׯ����F��8������M�})T��܎8G��	�����c�&?�V�_j�*����v`�,�O�kf���G��1iT^����N{7��`���h�$������>
`��R��!�p١�~IC7��F!(MƄk�i�����[��Z��~���v���U�,�%�o?
J����Dc��,��m��kM����CZr}��+g�zn�V���K���Wvר��x�Bt�p���f��"є$��(���<��h�I�qc �P�`�%�*�A5���_iw2��^����Iz,����&�_��e��^l$�r��>��2���P�q������	�~�BV|�z�`H^��%��z�tÏ����M<��K�Z,̤��ATW�z(�|��\��0"�i�}�P�׆%�៣_��aK10O�Rh�f��9���0O�D6��r?��P�OA���V[ަ}j��ҏ��ۙRj����+L��.��w0?{���P��d� �=�� ��6�˔��#g^U+I[����� �o�6l�u6�U��z�3��c����i���J�2�EwW�g�lp���ba�\Y�l^8V��\�p�SF��kO�4�W���or��)y��u=.Σ�]��K�5r�{O��9f��ؠ������	"m�%�.)dK������Z��v��Y<��#�R�R� "�h��T�Bb��Uq�5��&��н��.���t_��A7������A#4:����h 	�ɷ
T�4�M���GȈ Z��TA�V���s~�.C�о��ԾR�9s�Sߞ�M�bz���K�����ç^���+:��Y��A�Ax�>7Kso�Żsp
�"t��YE�!�J,�(c��U�7�X�d��qm��byV^��Хvϊ��%F3�m�o��N��x@��=��E��r���\O���������p��Ǣ-���̴q���(I�v�Y��c��Q��U*%ҩ�t�֒�}�Su�{�Ե��υ:���9z8��0q���r��f#����3�w��Z��ul�J�HT�"L�'/Ĵ5����� ��k�⪭<��2��.i�Q�νBJ��'Q��������U룫R�������%�V{�^�H�L��W�^'	��}ڧ�ˊhR�"�n��Q�ޏo,� �j�������s�r�1oO�[�8v��;�7�l����L�ґ*�7z�������7��������l�+ڲ�Ǹ��;ÂΔa��|6�uL_�L��0�Qy��ȑ�E��+#�Q�M�Y�Ɯ�CJF�1�D�V��3�����y[S���;�]v��qpCO��D3��Kf�E��o(��uA&}�݌D��p�.��]l@�Fu��#��2;�*��I��ĳĢG�˪��݅-p�AT����mϜ}�Uu�|�A�A�n�_ob�!�{����E5-o�.O:��|k��Bs��V���*�:Ԁ�[�'q ^�ܙ,���U6īty�A=��)�X����|�}�OtJ>�b?��"����f�.��<)���5��NΝ=.� ���Q���+z'[s��qz��<����Xq�B΃SRd��7����i���
�ʪ��8P ���K��iw\��U	(��H�;�������kq&�5�(k��˫�B�U�||nƧ�qq	��)��I��.+�ʩ���Ī0�[��!�,�F�C��P;� �h�O6�7��=�w�2Kǳ����f��F�#�����q����+M���|ء���|�x8`O2`�%3 ��~T�|*re�3*���3u$Uϑ�Y��U�\��:̔� �k	��綈���8���x��O��'�s1�6��HGB���� �z���
��k�y���/��2�N�c���� ���X��=�ቢ��L5�捴�[��>$��F8�2��{F���=/	J�S����}2%f�i�����n�&ѥd� �G�ZL}�,)������Ol�~V��B��i�[��A���H�\h�xɖ��T�K1�=���c���4�s42\��|��,�Pһ���C�n(�!��e��'_}[((1��y")W/[L�ɐ�92����<��esfĈx
/��2����#S�i�o�	�T���:T��� ƫY��n�T�ן���5�0��S���,�\-�r����dD�.�s�w�Qo�z�ލ��;�C���w�3!N1�vx�f�ig���F��<5V��F��k��ɍ�)���~s�/�-�L��i,�=U-%�NF>����n���TԠ2ԉ��嶈
��Ih��Jq�ױ�O�6��qM�z�"����˽j���2L����n��ޟ�����/�3�"����k���M��ep`o�v+��x�=K���NJ
8'�5g�����h;��ÂѠ���X l��G%)�<>oaIӛQʗ{�㩔�V��#��i�8�<n����d����W� ��j��������+�����?�y��i�� �#��=琁+c��Π.vs �΁��p
/���^��4�����^����@�R��Ծ�hl������ؔ"�@���QS��e���kS�dSqH��fw��%�f �C���J��U�0-�}���T{��:��lY<?�C1�׹�o���h�|���E~��f����K{7���V7�,D���R8!ɔ�@`����ε;[%�2�2%;l>�Q �$T�>;��W4d\lo�;)Î!��K"eq�:��^���o4�����5��ҿt5t)��C��=��/7@����M[�2wR]�~ _�9�[��s1^��U8=�������N�n�IW$�!�����`�GH���Ym�W�p� =�OB-Am��=�j}�	
'DR�~���8�C�rpA�Z0�^m��xJ�z>���RvMM��(�zL�0UI�Í7}-z��C�ǁF�(j��N�i%˙����V5�6�G{����3�b�١0��0b=�j��F=
�7bdQec�$�pAǙ^k:��AT�=8��#���`yrwm�p�ߦ\��^�E��M~}u܉����XN�N��[W��N��Յ�j=i(f�0�i�k穸�[�l�i�9��2��Z��y���J֓G�!��|���8�{*R�=��`��D��t(k�N��|�VF	m�ېq�����/`܃�{��XQ����d�L,� ��"w�g���C5�JgR�0�)���]U���RF�E�з�g7��ڈ������{*��Ħ�#��[�V���3�e���T�.>���CU�����%�4�����J�g$�5�v�TdM��l�gF���J�I�].Ih��;v'SէsSQ��
�����ko���@vņ6�I��������&���<Wp��kB���9B�O.�	u9E��6�TY�З�^T@�Dp�SRE�p�?��J�,Ph��6e�A�G'*�ckPn�����Uخ#�[����qT��6N
؈����c��Ԏs�������{iC�#�JJ@ͬ~�?�&�l��Vm*)v�HJ}ܤʍ@�Ɂ�~�ϊq�D�j��vu�@3���f ��t,����Ȅ\�D�*�*�=*���m9�Tx�5{5 ���~��g�k*���ʧpX�����Q��N~�Ȁ\
��h�g�,�;3	Ѵ���z�Y%�l��X�H'�Д���*w����=��{-�����@^�d�z�_��N���;y<��74� zD-'P��Y��sʠ�a���&��3?�F̬
�qv�P�,+v�3���pn ;�X9}�?Mfd Ƹ�����'5��M�Qn�8U�(�A�M���=}�UirsL�ī�&O�����hn:6!�vX0(1�z�G��Z�A~���?6�ѵ�f }��"�/� J�BA5V��9e�/��XW��K�.� <{�:D_8 ��)�V��^�[^Aa���^t������Ik6��ȗq�P��߾H��� �(ഒ�&��'=�@<���c��!UE���ئ������4F8�Ο;�Y�D�J�͋�6W�_By��]	0'^�K��k_<ٍJs|�#,�d���g�~�%�����5ݓ�vАz�v��B����{��} �]Q�XCtp
T�27�n�a�x!w�θ����W}�.���k:���)�'��>���5 �:��j��&�� ��Gk�-&��ƓS��R�\[��̒"�օ���]�И���I��mY�+�Ƽ���W�t��8�%�"Y����(	��=2���u-�'~�$�t�E0F���xk�T
 ,о������oZ�)�`������V�^�ڣT3V�ƅv�		gu�� gg]�0TstCJB���\��,P�Z� t��U~�E�I�*�Jg��3�@���w��m�K��E^`���$��`�>���Fљ����f��Bt7�����>��E���a��ta+���Hf���7��0�Е&f�Q�W�bf2�#?MC�3X��~��3y*J�N�b�y�j���*��M��ܧ��Aب���a!���������a�Em�B�魊�;�~���Z�
.�t����K@'IGG!8�BE�$b�r�㛉h��`�OJ!����-���C]�Qc������f�w�S�p~Q� Ti����-���U�ǅi���1����ʡۻ�����.6��4)¬x*n2X}x>)8QS����%�� &��i�II6�_�Z ��F
)�{}��G�y�%��aQ���Z�J���� >�V�{N&C��� ξm����p�L�������� (���6�b�&s�~Q���]����4�і�a�5H��\ nM��2^��ş+�
�~�����S��9�� �ƿJ�\L���_4�u��[�۠p��G�ad�)&+���>Ѵ���B�/���'�vt�-"k���UӝO�j]�h��&�C���k�M�I;*��k`�Pw
�w����?=�W��5�Ϊ�8F}g���:���5������M�S���-Z�q6�.�]A����N�)C%�0ޛ?5��y�)��������b�E.�Zq@(ws?Lw�pN&m%���+`M� [غ���'y#B�(�V���n����f��fQ�;���;u*�Ț��������9/P����(�*�qI��Q�.	e�,+�?5z����N��-�����wh��&��6�K���0�̟����Z�3�Bwq���A^@+�P�P,J���F>U�[O)}A��4U7�x�9����I�������%,f��͹5�4�i**��'.�1
RY�(��y]��ޱJ���G���@�ޞ4~q(p�̇���FR�Q��e�U�$����U�PJ|f�e]�TVaO����C�	��ʭR��~t���]}��XK����i���Z�v����3�EF�d:���G]��@�jGYh��� k#{�����u6�������Ur��W$��6�I��1���|�v�r�u���������P'է5�����RE�/�.�a��^��D�������IБ��}�i�9�������o�W@9A}0�1]���
�.Ͱ$J��U���X�1�7��Q���y�c®��Kb֤��%�ky4�:7�Jm����%3k�XBqI���p��W�&lU��,�R����
Q�^43J��@l�՗��Bn?W����y�ycY�pUH󹠱�)9����m-aEoQ�<�����}�/�1��L��d>�+6/��b�Bw�$��k�,7ʀ��~�kW^��V}��ÿ�����MY���#%�%*�A��)���6c�o�I%rI9�]��5�� �%OAMՇ�pB��<I�Z���D�2���|�-犲�1�W��?�sCm]���aJ�x���<е��)��t��krq��\ũ,��MaDx�Lv�̘���Z ���?l.w:�yd�����Z� �l��g��_|ߎ�+

򹀒�Y�z�n}<��TΥK�SY|S�\��q��Ʉ��H��9�D�l��_�����e}��T/,��>��/�=;�����ת�=y9s��skV��m�y���K�oP-TeXkξ&�K<���2�տ��)��}`��sq�8�{P��ʢΠe;���FO?���[�j�DŹ�c璳����vYir4�e�S��vZ�1��VO3��f���w,⛡N���&�s��N(!�E���T��h�Qv��4y�y
.�iR��{�{������,pi�� ��j�L@�h`�4a:���j?��Ie�"(ye����ڼ�2~xo����Jљ�.}����
�OhU0�zl|sm0" �	��p��n�2�ə��*S���o��J��'>̀��[�9�v�0<�Z���Gx�5�|"L�?�>��|g�k�*�TR��w!Ӑ~Vp�n�����I��p�{���v`��&"��5A�{��=��T8/��;�/�P=�a���`>
'��d�;��qt6A�m^�(�������GRY^��|�m�u�s�D� �gLT�=jq��h9���<_Oe�Ч�=y��T�5�|Q��ٺh��":�]�<���Hڨ5 �����o
��� |�U�#(�X�>�����-?��i���S�@S�y��.M���S��"�y)"�:{���UT;m�x�!�Lu�֔q���TUT�K<f2I�%3�r	m��3�x-�Ȁn�����5���Ԝ������#�Bm����� �e�r0:6*�����eM��r<�X�W@0��$-�㋥ZT�����C��5�bZ�������ѿ��(��8�ST8��]Ե�:2BM�ɸi����Q�릒ڂ�R��7K�_�%��w�š�Kfނ���
��N��pL�]� ���w���B�Ԑ�82O����l�8�F�z�<F�s��|�EX��@g�������MT6�r�$���۩��bұ�
�]��QƮz�+�`o.������i�����^�O���O�|��!���f��I�^��B��oD���'��s�8���w+�v�3y~�����<6_Ǫ9Iz�8՞���wg�/��
U8����ʩ[��5k�E]F֝�lf��Ô#�5v��)�)D�p�b�〆���ɣ\�8{�9'�r*n�|?5er�{���8��O� ��E[�x�Fۏ�^^cZm�+�ŕ��W��!��I��� �׊5so���-����$T¾�y�]m�h@�xx�kt��TH+�,@.�>�pä��ހ���F.����핹����K�Nq��8=�h�I�	� ����3R��!��#�O����;$�n�N��#Ix�f{�"�u�'z��V"z��̊llV����z!�7O��)��4���zyi' Z�A�=�C����_�e?,�fN$���y�)�*F�������:�!n�'z$���x鎶�n��c1[7� �����+���ե�bО;�t��4@��kwC���	��{R�M�kK_N���?��L�s�m(xy��k�nገG��.�ݮג���8����h��B��~mS �����,�j�QD7�8��^O�zČ���ڍ�����h�Δ���#����8�	�N:M�q����J26��y}��@��*�R�*i[�o}<�ٟ��:��#n�J��5������J:�����Y]UaBD|����}�&.$)[����O��jEd^��x�Ha��AS��w�!r���:9���)C[��N�$�I�{�H<*���o���b�D}t2�d���T��Hq��_�C蠗�(B�Ƨ'	�g�\��ů��
G\�@����9��������7�k|�欢*/�]�~g��<�;��.�GѲ����[7�4�`)f��2lP�+/c�v�}w{F׵-��A�+j��(�y���F�e��6�:�,�5��S�bz#Ι������J�2;�y�8R���e�p�E�U�&.��Z�^��cJ�G��D�6H����/3
>աL�,�<�#\��9|��� �"�-��ۨ��)�rg��|��g�@���9�5�;��=+(2�׺�VDe��k��}�	\��Bâ��Y�?� �.5�z��~��T؝Ԧrih��(�oO�M�'A-�OK�q_yR����#+AW����T+l��Щ���Q"�J��<�`�R����x�L��Y��BD;�/V��5%���O���0m��YHh.IWH1e��.b����I2
!��;,���B����vo!�W1:���j%�Xeҍ�҈Ó\�-7Eg��L�Ϭ�T{�ڦ����� vh@į:����x���tXR�H}���/�&a�^�ϓ?�{���d�M:����S8�a���G߾�
�r�_�D��U�8�����K��|���e�ktKI9��&b�F=��5���x}�8@��������0I"�I|["�#Y̓G �z Xb�P;�kl�<Cj_��}T�V���D�nv����c�\zk��>�H=�������Ǖ:/Fl-�w�$��������0ަh1�e�E�"A����<� ���P��U��#�
}������}`B��1��2Y�b!�~+2q�Q$��S��֑�*=YJ��˛p��"�W?�~<v��9�����'c׿�==��C��]^oǶ�斀�H��j������-�NM� �-z�'R�4N���2u�&�%�o�=�*��dDb����0̵lZ��4�FM���R�u�k*����,���H��Z�i�%�i��]r�~��XR�.��x��<�i���ȃ*���x����O!������ n�%�VX�^�\8#l�lK�;���ؔ�ؑ��������d����](1��JM�HC���tQ���+m���s�*�Ow����DK^��{�$����(�ꈘQݵ?՗�s�C� h�;�U�<9q㝯ͱ��-�z��Mӫ0z\��J,���=��z!@�h��y:s��;�&���ap�|�N[�������U5����Ex\s4X�ܶ�Q���%n��4�Ъ�y28<�`i�}�V^��PS}��S��Fu��ԇ��gh.�w�������/��,s?cbNu�~S��O��w�،�z�"OXC���+9}��9�P�"q_	��}9�|�l>&I��^��C6;~H�
��;�D!d����Դs(�؞y;�.Ո��B�[K�ݵ-y������Or�ʗ�u�%��@QH�O���p���+��]���j���F(/���J��!h��$���X��U%�^�i+.aWP
��ȀY1�V���.�桻�$��	͞��h����?�ڃ���S�O�2`:Ct�I�>B�Jf" ��B]x�ه�7[��juwf4x�����4�b��sE/b�4X��|\�cJ��U�j��u�w��s�H�*�\���eV	\�&�n_� ���:�$�*������w��~R�)m��z��@���A�h��L��dy�vWK�u����KlW�>�|�d逇m��L�3����T�M8���zM���G�5�\�	��y.� ��쫪$�]��a�9-�A�'I8`Q;:��`��5��.{��:r��w�z�����E�O�L~���VL��҆R^
�s��ꉎ�4V�k�{���SfD_�T�a��$�P��g��9S�H�\�:ELFu�^��<�_3���̷�2Z������X��rHUr��U�����8�"��:���>3x�r�/�l����蔇oŅ�L�1�&�"wS�G��/�#���_G�)��7�s���rJ�P���'^o���I��[�>�3�I)�Ҕ$a���/뀚��lwD��T��cW���Xx���35x�;�|(�W�z����Ï�f����)�Ӕ��	��Y���Jw�C��׃N������T1͗�[QI%CP�=/�G�%�~�V����Ji�!�T��h�ǲ�@9�"���ca�jg��$}�M��,��{�������>��_���j�ͤ�)�"d�+gbk��HJu_��9.�1��b�b�������V�e�r���C5�ud��K<6"���& �)�������ԟw�
�X���Nj��cp
LP8�m�����j�K���7��ɳ�U1++�	NG"�o�F O���M������m�x��l��$V�{;-����[� :��ɚf���YB�`����
�\�R��֝rqyo��z�9��E�A���R���_�� �ˏ�ﻎ^�P�ꓒ﵏����ȃ�W��O/,��)�����N�)o��`���SB�gQǼ��!+%����(7s3� ,  A���4�j�q�MtdE4����y��b��QӰ�;�*�[A릺�f��v�C[8ﾱ�n�uI�i�*1|}Ӄ�=�l����}a&����&����L����R�š��bNJ�
��gMt��>�.)ka[>y�{gfb��D����>J$]�]����t��0S30[I�
-}�]�f�Cx�e������5��Z{��N|�?}����a�ׄ���4�Rw��5�����G���n�D�o�v�p���zф�h�#ֻ�Ӯ�Ĝ�T��������!��z�?�aG[pY,��hVZJf�yB���T�<AC(g'�(�R�
���l^�<Q)�"%��>��FN��W���%��K�";�WT��F! �_�+̞)��0�Q��L�$��&;K��h���[r/�Ay�Fnr�H/��.Nl��&ӑ5P�q\W�ȣp�J��!^PJs��o����{#����S�㲲���3mF�-�;�t.�kdWS���.2����������)e�iS=k]�1�c�n^�N�b$�qm����NEi;�^��y>�D[ԥ�ǿ���j[J9����	�<�%<Jb���O�`�y�W?�^�� *`	�?XӴV����g�1�5=����'����Ov�����u��Ղ����h��c<�K�40G�=��tjّ|B��jȹ���'2�]ifn��HE��u1�M��xv�:�l�S��½8vLt>�g�M�Ya]iE2�l�m��$Q�� x��ʾ�6E�������e.�h�JT���e�IVF��)��V���ڎ��F<u�w%��i��`���D?��!��BD;0_=�h��N�����;��`[�R٭r�s����gas�]α�Ŵ3uB��R�;��<4ZCxfq�ֈ�;�@�w��7���ګ��0��� �v������ ɐ����$dJת��� ��XE���j�w��6�YM
=Q�0h���C��Yc��Nύ���[��ħ�.k�L���O���Fk�E���?�Q5��H5�I<fu�~��Z���4#�M ��߫`�uv�G�PO�SE�2��r��is#��ۍd]�s�7߾�L�]1��q�#�=;B��C�MB��O��{T�s��9����ŭ�+-%:�ܩ���$zIi�]�[�2�b1��[�a�PX�Pg�f��I��9x���vR�f�ډA��f>�^���"b{x)=ih�扊KJs��֟�ąx`贀���	����=Xu�|^��P�<�l��蝘�q�ؘ9����"�|�Z�t���]�b$�%Q+�<�K���ڿ�������.-
B���>�5��.O�D��t`M�������N�^#l���:~N����%�_kjc0�m���k�#I���k���!�Z���uS��^�	��Y��͆�A�7��	��r#s��(�6���D��=^c뛚L��edS�C�?b� �H��́��-�WIg|��h��f�A�@8J�QJl���K.��D����F���V��g�T����<��x
=p��R�{���&?ӏ2��d����g�።������A{����@�W8yV ��� �?��kgv�5M�F�as�N �rc|r���.�W	�����#I��`)`���<�,U�/�v�=��"j�:i]gTZQ�W�܂Z��9�\��`�8L)�6(7�������O��cL��-�^űO�������� $&ȯY�X���� U�y��ā�"5�p�*�&)_C�f����{��#�w�F2����j�i���L/��$&3D_q�M������o���f�� |��(vtP;����*�����M�9�Nn�R_u!��I�H���0K�&�aPD�>E]�!��(w�jg��e���!�+�-�%2}8�Z�(�ʀPSK\���lt��J�:��[�#U��	`�?�X��m2uQ�;fY���Kب���n�����1���V���i	}��M|1�|����%�qV7��5��!���%m(�Sq�in��S���N��$��|�6x�ƺ�F�HZ����o�!�gި�������􄥦���*�Xu)�6���o�T]R<��A�1��m@|9	��rrѦ8��K�d�E��F��r��^��eO�j֬#��Ϧ�� �1\��rӑ܂���r�>뺏��a�ȁzR�RrK'�����/�t�lj��	-���U���ܷ��>!�B��y�[2�M��ڐ�.�G�����̓���8�6B�F���k5\�9:�ݼe�V膏���>�nN����h��u!��ad��$��y�]{^Y3N��/�%�t����_�$����up�O�-X�(m�c�@�*g��gXn�N㒪זoK�c�ATW�ҫYB���� _��	�#��Go)U���y����X�1_B��uq�S�=R/���eċ�:wԼy/��š��@�V�{�I�6�8ߌ�6n���s`$����}E���KyW�����W)S�h8����J���G/݈���:˖��`��G-Σ����CC�m&l�dp.t�2��gb�+�=��oF+��S�J��F���6[H���ޚ_�I��Cd2/�23��#p�W�,G��dW�}���y�u S����J([3q�ݹ�%u��2���O���M�a�~�xhD�uT[]��
4�fB����9Ͼp'�3������f_|���Q�Cq֏�a�]�A��	G$0�$@��Rkw���ձ/�p�����D�C��}�)=j񬗴��;5�#��DY��L���M�-�d�-Ѓ��xh��M|��ki:�V^���'��r�Ν]2SfV}��M�JY7�sN[��Ѻx�@"B_���<~�c�,�ު��`��*=�[�����oS���0�;X��m�^^�m1*��AF�)��"������ ��v���5�H��6L���Zc2')'~C��I�Cr˫p+�׌��Vɐ?����ֈ���K�z�>J�P�,+��ߒ�p�� ����J�u�W�A}ƃ��`#����j0����-�%�i=ҕ��N����Ή9��8����{�6f�RL���B��2=rc4�>�%7�&��b:�����%��Ӄ�&�ig�½ =�,
����Rɷ�n�G��R��:-Ӎ�A\3�l�M�@���+�#�La)���)�KǙ_�B	F�`���J���ǲHa7d��dؚW�S�J�2l�n�F�{v�W}������qD`�uu�YBܰ�w��L�6ܓSߢ4x>f�g4ʿ�4��E;��B@7Y*̩4�_���w����$e�`d���߽3(�O����b��?�ɺ����_lF����OLR�m�}YiҐZZ	��ۻ%���:^�bw$`��&{;5,���E��<�DԈ����i7�-eQɂ"�Փ�{7�3���Ϧv+/����eE�����[�EH�&�Q;ʹ��p� p��~� �E����[������O�}�Ɛ	<���e�.h���]n�u����+x<��lE	�NgG�3rG�~ݔ��]�O��7T�TChu�:~�-+b�,6�]��m��NyN�-'�{BQ��t�{O��";prV��	��'%�+��S4$�="u�m����鱠ޔo��#�V�x����t���8]g�]�*��j��XuT�-�c�E:r��G��'bKqP���Ԗ��s,��}�=|-�o���Y�]���TMaJ�:[�3��`�-=`� ���H5uB-�Κ��Ev�FB ����E���-	�i4���~����r���`KJSWu𡙂v����wz����b���X�}�����")���ۄ}�o��-�+�X�@����#$�d����桍����[��o��ސ����n��'A�\�c�|$3(����6��*gOw���e�2�슐j\4�:�,��y�qe��^�q�����l��{`�1�G�P��"��(��*�)PQ�тk	T4R��z�rMϘ�t��oȾ�;G�ft�9�l��'Ù�.4�ҡr"���Ot�^�#|%]�|�#c�a����|����6%9���(�Nb��=� �)E:�(g�2�G(_\\�i� ������mq?#h�� �M�eWQV��/�h2�m�ͮ
PH���M��),Ւ�z��	����xF��~��YNe��:*�-�x��k�,Ö킠j����e�n�Ź�τ�>њ��a[��K�S�[��ʐ�R��?���3�+&R���O� ݲ&��pY���p᝽��*ܡb�,MA����ְ��&/�7�<���X��ĉ�^F�R�̐����K�t'�|cE�^����߾ƠN�z�<�GŬ"I直�2�A�w%耀�z��O�*���A�>)�_�1�6��V����h�ɩ��I�6d%��im{9��@���W�K	�+V�f&<D
��K0	6"���o)I���3�L�Pt�2.�8�ۨ�0Ls^��n;�3n�<��V�.�wGظ�C<�~՝�1`�ULA=�E����0���xD�}�S�g�����1���m4J��W&'�DX!��ߢ�$�#���~���s�*߾P������ّM���d��J����f9�	3`��e�t��e��Ex��|t���������"���'�ئԮ!�n��W('�gDW��� �H(�4}�M�K	����e�"b/���O
�p��,�%�|����(ja-4#?�ek���}�le��t�_(�ɇ�`s��Ce��T:�x4�D{��T����2)�#�7��(ph�(u#��Tr��6���g�OL���n��P�y)%9��6����3윴y�.�,'|)�X̫�u���lZ�W�M?�
�iz�R	�5"	���9�w�[�S�b�������v+�j=F^������"�Ù�J�2���D�GՏv�qK*�7H� �����S�L���/"�p�x���ppY��A �92i�	.�&8�I�����.g~�$�
���Au��H�]�-Вs�����џM|�ζ1���ؾ����n�0���<��B��ư��M93�7�"R��ڝx�m�j٩+����!:�Mݼxs"�%2>x��-�_W�LZ^�J��w�eԝ�ȕ�y����,uSbP�(��3r�:�=1p��ѓ��(�8�r�ֺ��n�/�89�es�8��"���=  �e���YK3 ��]Ί�֗a=�K"��vˤ�2� }q[vJI�5f�N��4p��0�0�դ&���UV4�C��Z�<���8�q��{O5�ݖD
��ڊ�+��S�h���}��������l���}�Y��q�Up�%R4��W&�.#�'!�`�N��z٫<2��֒�|d(�X@��3��H��j�vs�Ŝ�̕�bì8P�l�/��5!CH6B��&c4�	G�
�;^8��1PT����==A���l�=�1���eK���K�j��v?�bJ�C�0o��6���q���pS!_�24������H(�ٌ3,"�mI�S�L�W�,q$W�с��]�;B�e�_kNԨ��J\�뤂1��M�N[�	�:��+9�׮cd���`+חǲ���ͱ�끈�;��U��ZW.d>b!z����	�}�~ҽa�h�s�,���"��ͧ����a0F�<��ݴ�ϭ����D��e�jã�ԥ�O-4:�Q	����J��T\9�)p����Ϥr����T(�S���/�V@�!+����O�|m[�	EG��)Sa�|���L�L�E�ӡ((�G�ʞS�Ŕn�@�I0/3sC2�D8�ҩ\���n��^����H̖ޞ�9��(��ܯ��8N��K�0���#l$4kD�E�lh�-���F�p4- y3c��������1"�I��+�ԝ��\rK{q's �4�L���c!M����$�:����BNK�~@Q�LJ��t��|�Ba#���������8ҿ	X Oq�U^p�����xQO�2���?����OR�d���[��ⵣ�9�ϖ�*�U.��$�W��j>FP}9�����8&{���l��0�ͬ44���FӔ�?��\��U�
s�yj@~�~"�P��Bң��[@2Mԟ�C�h8"lB�(0���{v���g��JSOk��X��Ӕ惖Y��''�Mn����� Km �>tOr�n^�*�fX�.k�ɍo�2�yk赞�f
�H�#;b�׉h���t�W��	y��T�tp�@(GL];V7�����2���M5v����WG\i6ZG��S�n����M�Ay2�בdl�ȍP{<�F(v�pvt+��c�y���T�v~�I�.�7y`mE�\�;�-�$f�����'�#�� p��Y���t�K�7T�d�����
�Z�n�怽��"���[�fpgf\���s�a.�+N`�ŕ'݆~ԍ�(��Kc�'�vp�jWFݿ��µ�_��kmMWϙ�{Zgc����/��8��NJ.��!�}v��ؒJ�Y��Pf�uBvt�'R['o�6uy�8~gO����[����.�*f�&t_��rC�ƌ��h��P�|U盁�V�Z��]���-��秅o��t�������]>���-Np�h�������^�*��z�c���v*�3�1�W=���mM���V!T+/>I#p�U��z~"S����~h�-��s��!�>��8��I!�r�7��c������R"J`ӳ�2�j0��Y�����/�*'!�Qm_f��-�k� ��~������&H��gn���CqU >\��G�u��0ς���=Ufp���i�Ϡk<�oU`�����O�u��\i�"�+�wH+�'1��S�P)(�`413�YB�ăDn�OQ=�	��{�R���k'�P��O�2 T���}r���]�E�luI��G����8�Y�T7�<����JU,8�Tvm�!�a��K|�vVmQ;@��b�/��q��#[����:&0f4����x�)o���p�>k(y�7�K��*�$"��˨u���^2"q��<plm��qu�TVW;cz���)@��x�����*3��po�pC.wV�����$P�r]ֿ����;g��H]�./Jn�K!Ya^���<��S5>�@�4�����	��>g�����慆�L��cr1��H���|�&MKZ�Z�]5At�jj��/�\Lh�E��������-�(A�����/y)�<t�7)�М~H\Rds��x��)o�Z`�Þ�4��38�M�╘�e��S+o�^�i!rf�Oa������h�p^P�>NtO�h�|׫�=���B'@�ӭ�Q+~#�[ >���1� �}־=�.�.��TfﰰqS�-f�7�W�W��}���@(:G�Klu\(!o�s�yH0[g�Bݩ���$4cD=���1^�b�����-c��Rv Q�U�����D���I��t�O��䫰PH�E<�>�*8.n���c0ވ����^�Цh��~���`y�]�n@�s$�$֦{������q��lr��a
t�UQ�uv��I�a�v9�T@��k�2�v^���
��=(gw��=��G��G�e�R�`�h�|�b�⾿�����UןY����U7J"�y�4@n:�I!nD��`�]���!It%�	�,G�X�����y��k��]�\��
�HOW���[9�ܩ��#\ʿ��}UA��$G	þhR�aRDvQ7��P������ݒ_�h�5i#�H~�����7rsi��S#Ѯ��g�D]%�%rù=2.�$�o}��gАKLH�Y9�C�aE�T�h՞�i�Y'��z&D���!cUn�=@����-�v
���<v/���*������>WlP>z*6���
��p|����f�}������r�,�@N���6�<�Ի0^����}S`{�����w˵���Q���T(E7ObϺ���Q`*-)�����Y�7C��,H��K����C�{�Qa��H00�H� Q5�:�-a���c��%�ۯ0Ԩz����Qi��x54�$�(�Z7����Z$�ƃ�Pe��Yɲ0"7i�A�_@���;_�K���� �G�$��l���kBј;�^i)L�2r���j�y�H�S8f$a�e�VO��9�9����h��U��� *�s��,־�}��Y���˻(ͱ(އ�%
	���H��4��}031�4@T���U"2g`�a��9<�6>����8j�U��u��ω@�%��]"�g�ȟB�����n�z�B	�7�!��b��}�
�K�<%�*���j�o�&�1h�2ϫ�j���ɇe�-:�<RD��ƽP�p��_b��XJ(?�)��Y������Ŵ�zFU�d{�2Cح�@� V^%\�Z�т&��֧�������>�A�ی3;�s�R+�ֲ���=:@��>L�=	�(62�6��$�A�s�}Wu�A�:뗏�|�	`�ح�no���^T����؎��o��b���x,��9����N$&�; -�����9-wP�����Qü��Е��rJi/
��B%A����d���&J]-CD�c���V�b��RG�6,����x&�2�$�'%^j��
�]ud��&��O�;�����]}v��y�F���T�9���@�CXA�4K{%#����A=_5,n�9���f��_�@jzRip`�߬Nğc�n��8T�]�,�h y?��w�Qe[�FK\�m�p�u�D��C����A�(���Ҏ�����?l�S垤�T�#���w��#;��#L�9�4�s��Y����%|���>WeA����up����ݛdGJz+��b=�(���*���Ճ������99h�����6$���uN�!���}0Y|J�-�t�oe&X��[�<�O
gm�1'��v�z���D��s�U���C�����ŵ^Nυ��Wü�R�y�r�V��Y�Q,Lլ�R̼�t��������"Q�^�{�_w�M��o�d��6���A�p�G��ڍv���IÕ��I�a�[c��שt�mj� BHQ {j⡱�f�W�|1/�aI�ui�kQ,�뀇�_g'�;ŦQ��Z͛d�\
ȧ�x[5evz��㽀�	Z����^��������T���jZ���#'��tg�7��.��T�Sv�o@�&!
���	�@����2x�3�� �!�q50��j{��8ɸI�a2ۥfK(�ELd�IV�R];������p�]������@���Er�:0=ъ���~%j��c�\Hb^bs�������0�?��S�c<����7E*�{�б�����8z�p��wi���O��~���_kxt�n!d�m��%E��>�ҿ1H
����K�
d��O�E��;�Lq��`[���ģ|jL)#�}�=���x0����N[�+����p���n��	4t�}�� W��YQ�KƴN8�L����8�P3�|�T�e����zB�Q�-U����z�6t�4�T^Խ�/�s!�DUR�$o�ئ��í��K�5��_�]_	F�K��g�.�'�����K�7��\_=�	E������3�� G;9nQ;H�`�	Hz�s]/�U�����Gv�>_�Cs4,�+��A'��$��afO yh�@$�<��Iղ�
��:F�W��))�%�V�r�pac�m���b��g�D��֮[��4�G��+?�*��KM^�9-E�%����Uo���n'�5c�F���ǫ�J1�"`�L�D���\���V2�t:�烕:���
�M������}�e�r�3�"���[�X��G��A2	��BڊML_��N�G7b��� �C�Z���ơOIռ����s��n��@�/�R)Y�#cr��F:����tЙ��`x��fW��k\X�W�|��-���+ (a�n��\2�i����+���u�/A��A��~_���>4�p��,#���-y��H���}F�Xt��!m�ݞj0���GY�ú���D�ʮﾜu8~�NQ��C���$/��eIG�	��p�ï)>R�����8�1?Euk�yjz�3<���ov���#.�l��0>Mv}^�$���}Ӧ;'�v�ȁ�~�n_V��  �����.��Wsu�B��gY�zO�yu�:�*�B�֚��XHA�{��sg�k�@q�޾����(2�+u6խ��X�l�ʳ�RbfH�#{i��mt�����u9f�01��k���|pfq����ne�ѵ�YJ�����_ý�y�Xݍa��(mi<��MS�%��w�].��~�]�Έ�,N㻾��p�/�Z�������eO��Z3�E�MYY�	7^���E2�8|ؔ���׃��T0�78%�Q��^������h,e�e�R���>a�gj�x0p_=��%�hr�9b�����K��o;M��g�4�7��^C֤ޮwz+/��f,
*��C�L*t�<������������Q�6-jk���ҫ�.n\�������ӣ{�Ox�0!7h1F ?��ܼ��������L[%t�ni![I��"� �ݜ*���:Ug1��q`�ja[�<y�v�����~u=��V+C�����&5�,R����Ϸ���*A�؅%m|�q/f�)�f_B	�άz�7*�U ^�ys�ŉ;U<.y*@ޙ�ɓ~����b��7ظ���n��������˥Wg��Sʔ��-�um,��E(	�F��dj��p��4�^��4>�_F�h�F<�!q(]��"��C�^��'���$ۛ����43%1���*���v(u�ȹ-�����^��O<Y◨�X��Hʏj�����&u+��Fݏ(y��o���û�x���O���<!W�SZӊ竵6�;핁����^�Q�֮�� H悦�����7�S�b�œZ�$�5��[�CB�����<���ò���Y_��)&��IX�;#�OB�)�H�9�y��� �z�(+d�+��[��g�窷�x�o���f��@7��x��9���
J]❖Èu���1D+�F�߿��1�F��F���[!C9�\L�|Bs������	=%sF�Q]z�"l�:�[�uC�t#�|1XI�U�ؐ��n�rC�7���.a�]����? �+��E�ż���W����gk�,�,:.y������xV5T~q��Oe�)�Mw�>`����8e0,��E���H��]��jv*ß�N+;��u}�B�x��ȼk�b{!�~5l`�=�a?ZE �ġ̲�E�Yd���i�J6��a���&�N8g��m�A���Ǣ�*zŁ�Ɏ�y&��H�����m:�}W�aS���r�j��te˼�����>6nF��1o��g�G2j"a���!a�4�{�"��R�Nz#����ӟ˼:~su��ܦ����~?���d�m^g�;Q
c�EY����]��3VY	��[�v�~�Ĥ�E��<4��_���!;.�lԯ
±��.���,1���K����2(U�����ro��3L%1����d��ҴQ���_\O@豤间C>hB�����biv{H���kWm^�<dN��ϼ�,��ଊ�B�@�Lw�f��x�|�DD�f>�V�����6�_+��骥A�f�gay�%n<��]��(��,!h�K��L,[��:����U�7��oƄ�s��c̩$�Ȩ'��X�3�d.����؟��w���l;5��~<�� ,������̽яќ;*CkT= �IX�v���"���7��� 5<gD���-�5�ݐ���i�y�Q��aa�5����aQ˷b�]� ���G�Q�u�JǇ�EM����!�tF���1�|����gp&H��o)Ԟ`�s �(�ۋ��򽠄��|/�R�Q𒱨<�3��m �TJK4�ޝ�nEd��N��L��S�a=��)m5k.L��P�b@�|�T�M�j����:���1U7�v�
Cx����T��i&���_��V@q"�g�D'�6Q�JIE/pM೎32��Q%15p?�Y��gm�V�M�Z���-5�f5^�����1?^�8� ��N� sI+�����K��'�&Q����n�{�A���bWN��a�VG�L��ܐ�}R]�w��#���1�%f����c�}�� W��W�$�T+I�i#
֧�ɪ4�z�c��RDL�Sޫ��8����B?L�[�9�y7�.�P��г|o���a#�Ȏxt�.AMƙ�
5���I�_簻 ���H�IZFΨ^z��C���v<����;j;QTt�Ȅiem�k���;�-+t޻����6�����ʿ��JGt�*aR��i�.�D�DB��uȰ��>�%���[����*�"�a�1*l۰�v�(��+zַ�c��Ȃ�DÃ�>@T��?�}[,��m���)/�(78��FwST��|ʄK݌����"��� 
,O0���%�-��VX�������{�'N}�\�	*�-]�'线'K�&��y��Z���+L��J�u�)4g�׶�DH���v��=?��M1�d|wo@�oĊ��~�=����'�1�@j_����W���%��~.�[��W>��C0$YS�nU�޲R�0��:<V�<,�h���3@fe`87��Y��&0�t�Nʙ�����2��xO�%e�Ey�q�����R�EppZ>CG5DQ��M5}Ӌh�X�70�"�c�l�g�d����5<�^E�?�^���W�Z�Z��D�}�jz��@w@�T�qD�`��'���`_Jic	{X���O4�|��`����&:h �?%>�����F�b
I���b~/3�4�� �}�Iwr��}^ Q.�{IJP,�Rv`n�6�v�w�E�&+Qe�+�06��!����3�;����J��q\p�;ȼF��g#�2��́�%�����w���%�3W��OO�F��g�"�U�Y]�7B${S�b���:3
>S8�%��j�6 ��4h}G4
c���\�)[�C)�-�,�%�t�8�̻2%�]"�7�x�4G�a1G��%>,�� @5w�D�'��`6��u�#L� xXX6?��ʞ�7�W��ڏ����Z}^��Zޔ�O���ZUV���Q�k��'���د}��~��jUk�WB�f��v����u>�6Lt˪Ǔ��l��G��w��Ͷ�}�K�v�F�s;��`N(����YJH���/�µ���.<�؝�SƋ��G���Ǆց���ފS�m�6��{��z��:�tk��/��Yc��C(���f�}��f�r�Ѱ	�:"BQ$"�(�g{���܂r��vK�m����\���}i�ǡrj�zʵ�������w�'�-#��U�<�Eb:�g�J�g�~h�m��Hx��+z)�ƀ]�qj��r'0AݏؚX��\�W���W�0ƥ��/نW^y��d�!!5��Z�'W��;�RQ���)"(̈́Z	�U �3m�Cv"(�g���#8jg�&a,^�V쁍π�C.<�������*S	nGRc���FR���$� ��g%�;�y��2M���(bM���?o�9:&�(k��}fQ��&�|7딨]~���3�;��uW���C�Fs{�8�~]ϒ�. O���z\�F�;�y��?���k/f��`T��a�ö�%��.�`�V*y�	�H~�N�F=B` {�ϱ�6�Ё��EC��*���V&c�F|�#Q��T�4
�P�*��y@�"�8�>���Q�A`D­���X��6�5���|v��*�����%�z`˾��G��>��VI�\d���V4���(V{�1)ϛi�&EO�\�$ɠ�0�r�[~��FN;^�F�s�"� �a���Ho4�=�ȝ�eb�[Ű�R�<Uvʳ���<�j-�������Uo�c�R��?�ZN��p�FS�'w��*�����ɇ�Ӑ�5�)�w��}��*����������?��:ݯ�[ט��&Z�Vf3>�G";�Ns�`�M�sUl?m���d!`R��Ա�<�ܮ����TY����o`�33����3�]O�8ɤ  V8*4��;����w�Dﴓ�Sgu����S�B����h?���*�6d���%+���* 7�It�(���_�b����\m
�k�]
�^�L�Mf�����Mg͌�O1&��M)��U�P�>
�����E����:��(�r[�Nf���Lbo>؛�R������ �T���˷N'�<hErL�j *�3��u9㿹0ڈ�%�}��ˎc%5�J�����;M��ԉYt'p�"ՠ؅�;K��!^��f9H���ɟ �|�R�͊�/����I*�$u�A4�χU��������k[���P���qXD�ⵃRU���D�4�|�s�C"׍(!��#���n�;T'{�miӖ	ob��1�����fg��?�(��M��k��>�`����dT��y�qQ�+K�wݘ�.��V�3^$��j�9.����QJ�L������YG>F�,�Jo�gФU��n��3pg\�rd������ȏ��1�{��U<�Hs���L�y���1�8'���$���:N �(���g	�Sw]�;񴐰���KuѺ��*`I��j杉��d�"�>m���/3��B(}�~����HД�$Z�`�Y���k7��*���?�Inq�NH{t�Z�w(y�v�"o��ք����ؠ
p��.���T�خ�ՙ~��(O�U[��n�(���-��u`�r_�
a��@[� d��fZ���؂|?]�NN��1;��\��ȷA�i��!�K�U.8��ys<Թ�HxވC��!�:kL��[ЁT��Q¾F?q8�bI�.qQ�t�'FToU��4�~��|SI�,O�<Ɛ:�ԁ�Ԍ�Bj�^��� �#������Y̥ǢՁ 7��* �f[J�����m��q2e�誉�T6��$�'^����u>Ff�d!dt�3&W���s}�!��������s��$fE���'BUg�)��R#R�*�à��\qߋ��/:��࣋8Z`�p��8��;�:c,Aǅ$\������^�*!L��9Ǔn�P����KvZn�J%�������BdE�ġұں�W&#�/�=d i�L��3v_Z�����`X���*�Ny��8JW��v�������q�k������;G.�U�k�c80wǟ6���.w��&Q�z��?p[�-gL�i�x�9\`�%O�(����[m>��9eYM�*y�89u�Ce��~/O(}Fwi��픝�s�z��6h ��Ƙ,w$IÝUA��@�1��sȉ���}���*� ���jV�I֬D��6"�� ;�'�Jx�V�G��ׅ2��ؼ�T)��g����E���
��׿|�� .<�r���'�Ock踣��;�1斊D0A,��MV]E��80:��tk�F�,�3 %�i!�|m_,(��.<�%V�M��jwil��8r䠪t�k�Ο$��߲B�A\��:\<4�CUP�/�tK9�7p���2�Rc�N�h=���y�G�Ix��MF?����7"�+S [�(�BV���g-�|%=�QWdT��x{�����9ū�J�h_��Ng�pAU���mP5���ϯ��o�m����r΀��T�M%_������߿�#R���|h�.��P~>���m��S8���	x�8
��+H�D��{xM&$����EUu�i���ji�'R ���#���W�1��˔�ɦ?L6����݇K��MV�f�\�?G�c�[z^��~&�`N���Z�@�-t
0.�,ʀ�ׅ���_�ba�N���"wG��ի�X%���D���fQGIAt|E,w
��˾�!��v�����&Z�|i�HU�Q�ov5:��bG���{L�bg�{�WW��e�FM����2��A/�����@��~Қ>�'��G]h�O�q�S+�S�3h�K���,B҈���L�� �K #���2��<�	�*Hs閒`�OY]*�'<� w���5��7��T�'��N[O��׬x߽��(����9:>��Hg�2}�TB\�ÞԬ{��n�/�]S���YlΝڤ����o��sԠ�� �����gֱ�L�J�2��FȽ��WgS���D��s����U���%���De���a���7C�|���9�5"�53��S���	�F�sC��%�Gv9�� ��T�[4�ބ�+��h�s��$?�9�g�Op�˩&�$_E��I����P�m^��Q�R(R��G�?��1U�:ߐ�<�!ˌ�	�YLʮg�¨��Tv�z�-����� �^�q� YH4`�{+����2Ǟn��/WK����TF�h�Մ�B���J��is�S���.c+;f����G�Q��Da;iKQ�g��Ѱo�q�Z]F�� ;��/��=�O�,FE���9��K������A��kjh��Y�]���<Lr��I�uq�T���x�ђ�j<"�H����h_紓e<�����Qx[(��0d�_@��EY�~�<�l���|K��
D�4���JD4��pp�*��Ʉ�}�_p�����k�6�ͨ�:
̪���qr-|Q qBbդʰ������:]�_c-�{_;�$q#7͸(v�U�:����'8�u_���:�G�l�������W�&�̽=�g L���Ϙ͐��o��]�SLVO�����5�HjP2�x�n�1"�!P��^C7Gd$��Itz#|) )������Aw?֞S�7v�@cv%�<�VI��������;�S�g�s�8�ȭ���F o�X֋�b��~�`�;��x7��/���=TO��]��O�Q�@)�H,���j�l�ǎ\��~[`��+�%C7%�i�g��|�v�s�U���
R$0��?3�=�l{Im��^�H�-u�B)�a廎�t��5���O�'��eAXD�����ؙܿHN��2ւ3�4�|=���:��_��i8�,pli�L1�a�M��QBF�a�+W_�u��3������Def���0��tu+�e�@��H��Ix|�T>�_��sI����8`�=�To6�87��'�R����g�ǡA���-M�@���~Cт���3��.�t:������M�m��`ѷ�d~����z�F�l��Nñ,�%��7>�"�)��N�S~K����Oy��x�F�{=���l{�V����z���.c�?\�4�Soߞ�gl�����3�g�K!��Me
�Z@e9pG8���O%��>@�#!�ϩ]0��99�FgqŭXZu�ECX_���:����V�Ab�����3�5ֵpT���v�U���� �u�cT8�aD]��nc�z.v!���g����˄���Zz_'u�;�?o�\z[?cre�7AʪG���G�Mױ�n��OL���83C��ڀ!yFw?d�#�B��]�3�J�U�XC�{��N;i�}�P��i#� �MD�8�Q#2�G��'��i�gv);T�*�����{O^�&���rD�z���.��(���sԨ6�h���ڀ�C9��\7|��͍I��*_>�vB��o:Z;�Q>{cv�K��bp*�)qv���eT�����4�{;`��ׇ����R���\/rL:Zc�)��Co�aOdX�Ѽ��dEd���"5Ҙ�%tI����0�[�ƅ`ÒݎJ�F�'jvw�h�Qo���Ԣ���5�dѩ�+),�y�"Y;#=��G�u��q9W,��j���y�I��	M�|�X����i�ke��VN��l�� �3M�2�y%A.C���߯�-l��lIA.
�Ȭ���< NظTL��{i�%�[����'h%��̇�˥N`d�l�51�Ϫ�br�ζ�b'H���>�D���CA 5��~5�]�ŉ���e̼s�{w����H�����o*��� �Ok�e�0:?�F�n��yD1�n��m�
S�>�q������D�]�@p��, �Z���h�7��g	�pP�/w#lF%��'�5��8�I�$������n4T�Pz�]X+x��\E���x̗	R�'@�������Ē@q�C���-[*(zo�6���p��"���{��U�.�
��e��\Yv�Xh �1`h`x�Q�.����'@�$���=��k~�p������딱j]nb9,��˧^��x��z��F~�:���ͭ9�A����NB�d���Ѷ�!�d��l!�a���>)���!���9��1>sUYS�nmj/��8s"v�M�]�f0�ƻ�w�q������_�J�cH�6�W��yM5�U��՟���F�זZ��ul���r�G�$X��}�*}��s� =�E���C�����K)��n��<��(�ը��	W�L5φ26������MMkxF���S rY�lk'ū@�I�����'�Jj��Im��gKڰ5�ʗ�V#�R�~	�7����!�N!?5-���˅���ڥ��������l;j3V�#R0�9+� +�i�
����Z*��ژ�̪#ɂV$=7I���O4]Ѷmܞ"��''��wiYN�w05ؚ]��C�'���OQQ+6+�?�DՖSu0-�W���6IgC����[Gy��^�Z���~L��΃��y���C<��������b���`�xw<�0o��+�@V���?�@�L�\������Fb���(n�C3��1�+���L�גZ�u`/Czjqkw�������܁�+Լ��T�� b�ڶ�	��N���{| 4����YI(Y� K��,z�S���L%� Ŵ�!��~W����,uz�3_5�O��.��bk�B-�t{�F 6�5�,b|���U4�a�Z�aF�^�xA�xn� 橪A5A i0��ʟ��*��\%��t%��2�AbR(�-����i��7 �w|~�=�1���0��>�?�{�q�,��g��W��j$��(զ��^ZQJ��?��h"�2D�9BP�V��\�Z�.��੩"��e���)K�5�w�X�����R����O�����K�H�!r�+�Q����)�'[��:�ҸXN����B�<�����YbvKXl�^�'���V��?�I�{
�ʶH�0{4��]��C�v�nV�p�Ԓ��w��)�P��UIgQW�Ҿ�f��}�G�:�!�,�J����0�Y��=�B\��b5`��5�7%kZ��:[{��J�ß�W	���cG����~1, ay��?y}%�v�e!?�Ȟ��F"nx_�w���S�)Y3�e�֍�>.>�ozĨ'��JY��&�g���@o���;Q�'�[9v�o�:9���M����|���Yr4�6;��>��e�辱垕�H�̄��m�,� ˆ�aa�Yu[w�hg���(�?I��	JCq�Y��9�G�f�Z��Ǒ��)�O��U����O~m��Xb�����y㍬�ϡp�tk��Ȼѫ�6<����G|�Y���2$ ���Jl��8�ؓғ�kZ^��X��Ɉ��A� �Ӫs� &M1v�÷�61Y�^�:�@v��� ~�rR����	W�jǙ+�+�=E�Kc���'UۈsG:��D��P9LbƩa}�`�k��s�ly�#w�X��Mz��X�(g��]Ø��[G����
��TЖV�x������P���v��2��
�?ҷ��	������6"àJK�u������y�B?�95�Wh��8��w,�U9ɘ,�c�7)i�A��pΤ�+����P�ʱ:bP����e+��KȢ����6e���pE�A��VA��*�(Lpa(�e_6������Q��IeasZ��N����N% -ɥy���u�r�@�4=�7о��X�aM��(�|���(m�o�]N`̸���y{�K�裘�3̢�I)p<��=�j��m^�*�������	M*о��Ĝiik�,fltr�W�����3���$�uy:V�B�[4��F�"P��mo��X���R�W��t&-D�f�=�U�tmv<@������<��x��d����ӛ�;�A�S��w�A�P�#�+էN��
B�Y�ʘju4���d�D߉��#�0�U�*P��n���s��~5�ܔ�Q�9�+��?c�8:�\�Uȡ!Ϫ������ώi�������K:³���G;��\��H����r���ͮ�x��҆ӡ����wn� ��wCX<��G`.O 7R�z�3c�S���,�S;ѷK�O�u�tWPp�T*ɭ�\'��t�d�W�K��DvDJ$={]J�"
ƴ�`>9P�?l+��a
��5���%p��IkI����_�L�ж��v'�Ƕ ����B��&��`�Q��ߵ?��m�ũϐp�~�&���Q�L)Sez�?�ߎ-�}�Wlqeg������S���-��E6!L�w�6���Y�0�D9h�^�4_�v�T���I���ī�
�v��ϲ�E���W��o~9���~��L�\l� ب㿇V��7��Ec	>\OX�jJ�(�5w.)�)2�>���y��X��4d�X�i����Sg�M���U�)"����:�[b޶I�[����Af�A+��/���݁o��d�� q�bn�$�߳��/�v\_G3<��7�tP 9�tDήr�ߴQ��:˚�]���}u�P�߲R����5h�����>�-�TP�H��v�s�8���f�^,ܯ��	�g߼A��Ip��a�F�G�	���4/-��gE &��BYN�]5�
�I��J�*h�SX�g��5V�� ܃�_�����ٳ�u��V:��f2�[:��z�p��,x��]��}-f�%6_��0B^��8O��jS��0�{`qwYxk�Y�59N,�}m���,�Q���;�b@�#��wq&�07�$.��#��ׁ�4D:��N���k1΍\��Lg�A���!Di�>]��M���g�
�wF���^�Hj��
��e�k�O{���<c��E��~%[�T���4u�C�Ӥ�/�hr�lɞm*,�4�T����;~`(0zx�GQ �D�5��$�V�5�.�f88�8';.\t��q�q�]�Ef���{���D����E���ǯw��h�^a�F컪j��><�I~�AS8KcxN_��v�a�!�Tf�s���BB�������H ��<nA[\�b����l�y�������V�u�bح5Y:5LC��*��;�0�:��g�N��y�2N��O<�ҥQ�
�3�܄žU$={����(Q Z̦��K���B5�*�o�e�O���$�/*-��$r���G��}����B���,��ύ�	A��p\�S�I�$�|���v5�r��\����`�����INju��*��"\ҟLD{)�����f3A�JQ�U[&I/�x�9�h]�|ó0��k�?�pM� o��q����D���@m}����5Ճ;�8+�{{'V$[}e?�+c�����	i%2��aj���"f��$��އzX�X��dd�:�q"m��8�q67�˻�sݣQ'���V4;��Q���6e?��:��p��s �Q7iԙ<1�+_�x�8Gk��,WfK.�i�wl5��9��g~(;AKyg�|c�ir��A�e6�h�*i����!!%(	�9U�h���<��% ;�7xBW�-�3��.�@Q���~\K�!l�R>wۓ�[h��s�����mT�����_���r�gb`p^�^z��/�5 ?6	�9M����x�?k�I�k?�ʅ���P�;,�	ʂ)�����k۵�w8!Yޫ�5L�Y�瘨e�Y�K��hk�@l淆�˫K�����?��+�2��[�q��]_uCʀ�_u�s�jD��V��snݛ����i��ois��C�6�)H�]z�����ꗙ�8��KCCO\2�Uz���ԝ3�ٚH�r�X&�*f����{��Rl�-�@��b��IS"��`Qf>�B,L-��齓��yu����ڲH�����' 4���#�b�w	���_A�����DNH��s{��;YT)Ea!����O-��9��E�i2��D#��|�B��z�f�f�~{���y�	�eVyjh�,w��<T��H*b�~���0٘V��8�N.��Ժe��\B������̙^�R��J�=�h��>���C��'L�����NVO���E��x�R�:�S$�y��ӹ"����:��aV[��a�3����jm�=�"~ѐ1yX��!��'BE���Vm%6�ǁ,/��~*/�Q�����l����6�S��A�aӘ�2u��Z䆾�)�Ď��C�=9ߕP�<��>��﫪x�O��	��^��S�� w��t잧Q��|6�����|���!B��Թ��MB��XD��dbaS��W��+�$��z��M�?�I��6)�6�J��8l�6����
�< ���ӿ���g�326���~�D�3s�^��Hz����<?�'� V���3�'D���4[���Y	i�A���AK���0���]�r�����P�fX�ÿNT��D-�e4��V[-��j2�Z����P��{�j�!�!���f~ڸ`�����`cE����Xԯ��Q#�~gq�:��X�V;^ֺ�OKC�]6VY���A�����uYVX�e�&�G�c�	�~W�a�,`0�7Ď%���QRU�#�4�V���u�QF�h�����5}*qpa�2��7�zZr2a��&X��;,QK嫡�����	�'(����o[
��j�	g�,�m�`(����VyQ���D��e��F��CȎB���g��R^F{A���^�Djѓ߆U���Q�:�jui���`���(�K+GѪ2�&p ����f�-��o�t^z��"$��UU�slv9����sC��d��į�Y��C��oG���ĸ�|C.ޠl�u��s��JK��E]�EO�=f+~[�܌�rl�3BF�"
�v&�ՔT�dF�!��|�U2ǅ G�f��r/u�s.��=����4pW�3+k
������f�㥦��^��ßBΒ�l_�����qL��Ko�"r% �%8v�p�����T]#�stܴ���y��d��G�67v�|[��7U����1��0��s�N{��)��"��Wn��`�5�=�����KH��k���[j�T����_�-�Ok���
c^P`�l���h
�=�F�s_ρ�V����5�j����x�P����ru_����d!��O9̃��<аzH�l�ʢ�i��?(��Oi��r�.���S3���ڪ��6�#bx�yP3z�塽(#ѧ�6��{�4Bk�7*j��9�Ile��iG���P�˼Y\�J�IR�ɫƼ_9�!X*�r�����6g������=�-$Y��Ҍ�N����\���������֏�o1O<z?��\��9|Y�a��R�z�m�uʬ��u��0OF��'sgm� ��V+aek��
x�T�[�ca���8M��8>AOol�#aK(�U��=W��� �3k@z�;e?�gy�G6q-�"z���o]F��fֆQ���6����;�4�W�$kn�D}�#�n�����poň�<�e1�ޤ�y���|3Ժǔs�+�(�0��8M%�t���%�p]��}1T(>�!}��708/P����P����jA��RS5S3�aW&m�=K=��2G�;l�e����g�R�.�Mp��+�>(�1j2g�c9BeM�l*�*���B��Ff��c��E`#N�}+�DҲ~�Md�t�pR�TRRX���!H��],�n�0�(]����yW���f�:`M���&#��]��/�	@�_�P	Ϥ�d���5#� �8<B�\H��G��ۗRAⶳ}�3��w �\����,<>��v�9u����f9"��P�O�o�-_���/h���.�ӓT7�N�IZr'L�5ىG�4==�������5�����tj���)��l�3t|qV��i.�����z(�}�$�Z��m�qT2և]s�O#Dc�Y4�7�y��wH� l����YI2��p�I�(�U�S�YI_7����,��Z)��[�Z굌��QJ��]?��r�,YY�`Y�ֿ�Vp��[m���w�Dd���j�%����I�jx�n��P��*�H"��+�MT�����:�۲�����Ɯ#��j���xx,��}Ǐ%~M��UxUr/���ղ��#�@y]-��"���H�<g�҆�ѳ��ڲhy��	�Hz(��q������}J�NU6�����IT���^��n*�i!�mJ���$:F%�@����G:
���E��"��OlDY��T�8�U殮b���u<et��<�l
�n3\�!pJ�g��x�ȱl�8�����kc�'\9��!�GKS��~/����P�R����\���Z&��/���5��3�-��e	���	*�&��W�+����b�,k�aw� q�[�R��Ư:����$%��z��hY*��ok7<�c�@%�f2��^7[���/�NG;�7��0���1"��V޹/�ΦHm�T,�3g��0Gw�?�p&���?��*����2���� �+�VIτ�Bʿ�{5^�1�����
�����5�`�߳�f��+)窑B����kN�a�"��(���l�JE(4�������_ޝ�b|�tn������3+�F�E_���Ɛ؁ �G���Ϲ�/��q^�&U�Е���c��ܢǺ�]L@A���ˮӀ�γ3�R���k��b���c�yim/�<��a�:#G��0�YjT�p�������F����q�	-�i�ޏ2��P�t>��Lm`���v���R5`66���{?o���+�ػ��Ƅd�1O�m����N��M�P�/DU0f����}���suQi�M�[m��7��|���!��ȯ�d	�MQ�Bb/��h��)Y�Nܦ�fM�{��ߪq���	Tc�/�0�̭��,�L{lO�*��^�Wʍ�=s�7u[��&=����8��Ϸ!Q���rHilw��H#�w�0����O[�N�T���OQ5=\ap��ҏ	r�oT��l���;�<��R�HzR6�ΰ�d�qBj�Zի'�-:4�:����T�ٟmX���3�-z�ҥ�����t<eT)s��87��eϯM��e�kt
����d�u�Eo)�)fkԶ|3S���+�e��2����k��f����Y�U �����^ ��n�7�/CXl��TpN����Û=��9!|�3�Gh\NF�]y�6��N�Ի�)����sn�9G�a�|�9�C�G� ���s6��<y�׮4G�M��$	p���0
]�m��9����~N��Wp+P���̇:ɝ�$So'�Ѝf��
T�4�W���]\���|�2��.&��Eo3Ԝ���p{�e�_�� �l�< ;~��}U0��`q$D��U�ʎ߸��v�ȯ��V�J�4eH�g���i����o2����mo痔;�5o=n��`�.���Y=�d-NxLΠ�ͦ��y~�t:�O�K�yԵ��YXN�`"�x@M>��b[P�պ�(&W�����(���
p4���s��@�z��2<Tr1I1�x�uԌ<��%���F�la��u�|\�����[%���?E ��EG��I+:���[Pм,<26��x{ق�|�� ٜ�{��9��֮ﮑ�Jh7�*8�qu��	Xe�pkdߑ��[H�F֌9�~�F�T23f��D �[4<������~{uA%.�7[�������q�xc��A6W�
��9ka"��F	W@	��h�=Pw�������u�Q:���C���H��*`9C m���i�X��q�2�_�����*�Z�Tn��%�h�@��q� ���>��S�e��d
8sի:Q�S��g��R��F(t�@y��H�7�>�o���G���nab?��c�\Ya!���k��#�AD1�s�A�u�~�����p'rl$���9G��N���5�O�W�fp��n�/q,��w��B��[KՂ�Z¡ f����̃ �(IuИ���DL�vF�TO��C~z�����c����� �5=���rL[�q���[P0�w]��t�$��鍹7��*yWxTk��H*��Q��55���ˡR&��|@��r߈5�]�����L@����z�LQ$�t��ۉb���#7����sr���=��uN���S8��S����v�q�1)��ٚg���~�y�X�) c��C6�P�[NP&�_��_J�ԥ�w�-`���^~B�@�w�xg��ٿa
���6h���нk�D����9��7"�u��c�����Z��ܾ���ƕ�}R��Ҵ.�56��xI��-�k�,L����a��o@������r�`��
��"��	f*>
��ȆO흿��i���Ո۴�C:!r!)�s�V�-D��H��9�<e�:8��y���AO�	8��F���m�p7\:�r'��8G�]bp̖3:��@Ұ�՚�k��)f�����Q��f��nH?�,��[~�T���Eo�o�}�ɔ������##���^�������E\���ʼ]���_��;~d6>�� N�����"o@���R,ZFq�S�������Ly��QC��q���rn̒`K��,Q�o�4*���չ�V�!R)�U�B��[�B����/D�`�� U/A��ڜM?��he1�R��ǐ���-�A��9��&U� �Q�-��6V4���S�����m�aa�ǔ�?_�ޑ{�?�y~	bB�S84*f�*tss(hsu�\���
k��f��
��icqq4m������;��4[}^���-?�µ`!{5��]|�
,�>y���9c�����R���?�O��͉OZ�o �2�.�<x��N�+�oZ�Qa�㏔�Sz�DpBy`��x��޼K��Ӄ���F���.m��Q\��O�öl�����·5�g����绐�{rL���\��Y
�ڍ��f��c��S4�$#�@<�buO&�،SS��w�!������XO;�4��t���#C귶�����b��[�^��f�KJ;h�|}����QLHET�Ǻ�ql}�v�z ,7��W��.��*	[�L1�#n��d�L|*�V݃�:�W-�ʓ�DPP�����O"��e��%uH���&爙Du��uc���C�c���n׀�ݑp �O��c�����e2�ִ�j�v����%i%�&��Jɶ�}��D��J�8�?�ɢd��(��E���R%4i~+�^k��-�OQ.]�ˁ�ɭ���Z�D�7_T�=���S+<���.�|������V�d�B��ø�49,��E�aH��gVweR�Qs���GVw5�v�����ۜڻIF��H��k�)z�p�����]������1[�m�F�����^;��R�%f��x�
�k�����ӕ�3�\��6�#�Z�c#�H�y��yă�ڰd� ]�}�Y�aZ�O��b��wؘ�--��.�%�|����$AU��ﴽN���g�zK�4΃r>.����Q	�qbje�ON[?1��c�wDL
��Px&]�A�̒��p6��O-�nac���k[["�B'V�s�@�ɘo�5�����5�%_��ۜK��~ɴ���[�ھ�����	8YY�G+[��]���+n
2ys���������S��J���,��K2)�p�P$*�*7/��	H�<$A�51���1x�}7�s�C@��g�I�$�/P�/t�zwr��<
Q�u����V��K�*G$ؘob������w�?����I�$�TEs��?Q���G0����u���W�("$��`��U��) Mg\yX�Cx��l*����@����W�7H��-�^K,�wQ����p��Ο��#��R�Q�	����jBG��g���7��[CD#N�[�Y�߈��W� k5٫Ъ���D�k�zx��Qu�ٯ�P���� M	\�}�d.^}�Cv;eu��6�H�X>��H�vn��c l�P�N��:��">��'�͏yT���G���a����z5�\�7̅��+%��z����w� �GG�&��"��o��`Y�5(\l��n�ѡ�P�B.�]���ɶ�
��?,����Z'���T��L�%^�W��L�a��e������ri3ZD���e���>�����i�L������n�RO ���1Nf	;��	��55���qҮ���H�o�*C�4o�wLz9/�=��-^.���h����^��U�'�<��*���t�D� D����`�h��p�X��D���,B�l��:�����ʾ��ͨV�s��BF�3�"I��O06a0W�Ar�1��d��e�  zKZ���ŭ/��I�W�è��F46�9�'v���|H�^&�`+@j�o��
��wS��K05�#�_c�qt�zb[��}7�H񺒈��m�)1�ilmt! j9��-��_-�-���4E<R��G;�������S.��g��Қ�孲e��$|F���|��Hۈ.��^w0*61�Lʶש$){qX���ER=�g3@�ny�˘"γ�e����B?In&�?��F|fb�R�e]FwF	X�0�)��kK��gީЂ��Jq��đ�����Ră; is;s;�Ĺp��5�K�5v,J�6��)�Pm���4�VQ�x�����h��{�U7 �#�Ѩ^Pq+����!C�ζ׏}~A�B%��0�+3�.=��U7#J��=C�)�O�V.�����r�=o��!��XŌf���﫶}M�"�4T&㰨��#/��M�{RsY�Τ�TV����ѣL�n���[1*�5�~�(��1�Ϭ� ��F�� �O���&��������hx��!�r��B�b�ٙ�cС+rn�"���G�������rN����E��HE�OwD�,�qS �q��V�K(��}��o���~zH�L�Pq8^u�	O�ԙ���k�'�y퓲���Wt�/p��)y�s��g�EU����lK8i�3���"qdKF��R~�Bz�7��2�y����#��`zi�$=r(���#U�jr}�����;����)���tc
R�Eu�;I���'��ܕ!���V������n��p���H0h������g'�B躆�<����R��UR��<�pѾ�̀O#y9����[�F9�����R͊kV�ר�~!�c8�X}���y�R9�� �ý�%��J�Y��{A���(�s���#����%CC �~�!��\0E��ݦ%'������\�]�����HO�f#�N'{����W�, �sW��V��bn�(�t&��Q�a�7�Ӕ19�/����l&w�J%<(���]��eSS��cH��Κ٧�;�B$҄f�|����⁠@Y�#����[��8�)���
L�8F�X����^{����$sR;����><��.Vⰵ$H8�4:���-z��0����T��DS�lS�\x�V`b��b�����
v�T*�w �� �#X�����-�bH=���{Ֆ�+��(��t��R�i��5Pʪ>�B�AMFm�K+��(�E���9�u�1����܀f�DYD^��a��Y���m��I��4�RHt���N?�Jm>>�B�fM����`)9��y��@�h�S3���c ��/#Mf0D�lq�kMN�|���5�h��l� H\S�Ʃq�F�᷹�l�9d�'s�3�&�����c��ad(�1���l*L�U�K|"QX؂Kk�M\�޻z!�B��)�'�T�����2���a����P7֟��:����Y���7� �k{�ӅƳ��+O%�\S���ca�<sA�O4`�x� 8�ӑFd�q�4���%f�rޮ�����Sė�g��&迦XM��mJ a�ǨQ'����[s�\�cwd�NT�ݖ�<f���{�a�H��ǵ��f�f.�J�N��+S�N�bG$�t����X���j旚��1�>��2��'�X^՗��vp���
ƌ<�0��0������	"C�2��O���l\\r��� ���?t�!�������<YzI�H�g��T�^=���3���*�d�\&��p��9�N�Rj!��袑7S�&�s�t���<|��y=��W�ME-.XP½�����,��g:"[����W�T2%.�@��Oy�@����:�֥�^�N���Z�|�N�L�.��ul(J�N�������G-=��O�@Ʊ�����^�L�3\Q��pymeR]�3�a���%�����:w�#+c�M^�$xD�Vԣ'��;I��t�"��������T�*��y�%��T
&Ԓ�US�3s4!1��iT<4"䝀�=;"��+�MB�O��C
����
ҝ��_K�[KE�OF�B�~DV���pl]j�EF�9{HZL���G%�l� f�5h���IP!��#d@��u{�u���	�+ع3*t⵼,
co�j���̢Ǖ"�-�&��4&�ʗ�=� �A��-��~�ro�����'>�����ۿ)T�m���F�zg�R
��hz�̖٧,2�=��0Ѹo��m��M5��~�3��� ��25懹�=��ed�`M����K֮'�;y���0
�5h�� 7<�a�=�}u@WY$�9D������)2�0�!Gp���JUj�!Bi7D�+�Xpk���z����m�USՊ����f%��䜼�/F�Q$���Z@��ͣ� ������ 9��vd#��aEMq�2� ��K6Q�O;�*��ǁeE��Q�+������/�-k���1��ҽſ��#��rS\�7�ؿ8P�Tt ����	����IcO0����9v�%X|C�0 �' ��O7�q{��Ffcek��	$���i-`��ϛR�i��BɷG�&)]{dT���8qm6��|�����|�X�TFp�ݏ���Q�O0|����6Z�S
����
u{W�ƅT����yɍ������Q�J�4�G�1�yڕ롫�N��� =��ԏ`\�+r�U��%9T�q��0����UtpP�$F���)�1�:)�'�/�m���x����B�`���)/�r+U��5�W��IB�أ��FX�I}�0��b��g�0���"f��#�IL�,�J�e�2��qł��Y+ܼ���r����1�4s�pK�I��m��7쟨���W�;]�X���-�����E^�U<�{ѵ�	l$�"#Jި���ʚ��!�6�F@HY�E�+�������_?��Y(,Cȑo��d8�8�%�H\���9,�a9������arד��p�#]0�;��3H&>&�E��]�L\�Xu��$v�E�I5n�㞋�,�F������
����R�s��K�Ū�u��
���}u��\�D��-��2����hJ=���Sٽ�SJ�ht���fZ�ԂXp}�B8m���x�	�-�$/:!��V��^�3�cv��5��X-��:�Z1Q�WN'�0��σ|���jn)W7��P���fo��*���F�aCVD���j�����l)4���4�Ջ��=��NT�{��1F�H��W��m�x�b����Xt{����6߃޸��T�x*_�0�g�?^��  �&�]��G��i�_U0$݈:H�mY��%�TrYd:ho�/�6L�����&�������^���&�~c��%��Z#�ݵOBթ��i���Kd3��W��p19����L��ȰR��C ]���ylj��P���5HP��׽Z>�ڍm�e��7��v!��I��ʮ"���9��C�vY̪ZD�ƌֈ�@�1~J��옟!A�af���]޶���t˶��ҷ����0�VUc��!?+k��qO=*d���u��U����2���\�-m���k>��g���ݼ,[;
Joݟ��N�S���(L�����E�k�6]���:���BS��"uֺ��n�8��A�����ڏ�`@qS�U�gV�1������4����S�kx�8���X�=ntn{�K�R�H�ձ[q��
���a�Ɓ�P�,L6��%U��c������� @������E��J�iڒ��@W|[z�h���\'��N|�- 
�у�R=�3E�e��F����xe���]Y�G���Z��%�gL�0�)�܊a9��A�21�E'Y���{E��÷=B6Y�E� ��A�m�w�F�ɏ���v���5!�3�*v�������R�����a�P��
�R�w�0�� �t�	
ZgJ$��Ύ�0�ٍ�P_��4��w�9�K 	m��K&܆�����hNq�V1s��{Hr��plH0E���N�`��"��M�Le@�w�G�b][����7(�W�̻c�	�bS (�=�-�>��Y��q�윜l ۄ ��)i-�=���1����0����$Z ��9����l��n�z�&��? ��� ��4Z9x����}1N��}��ף���]�V����q5�Ѕ��D���V��l�1���n�L0te�N&�>t�{vnCO{Ԗ� ~��+`�pͱ�y�m��������E���Ab As�9�J�I�"1��+g�(g?�i|�8_rB�Aei��d"I����G��f�/^}`_3>�2���������Ϡ���E�@��O�̫j������6Q��l�_�;�(p����h��G���c�Y����&������P�Y{��~W���{��5�[����3Ɇ���>C~�iFf{G�e~�e�@`�d!F)�\Ƽ!%'�O$B1��	��Z_6g��|=h@I���hK��I'+���'$8����qڦ�N�Hb5�!�'� *������^�ĩ7:��jۋ|�އ>@��")��B�Ñ6l�T/�#{.�T�1t2<���K�ˢ�Ⱥ �-���t� ���Ϊ4���ܗ[4R���f�`��d��x�j���-�8��y��$
9-T�K,Ԏ�|��{d�������w�3�3S�k�+���f�9`j�����~�|���KL/f�K,��v>Cs���?�blu��]]t�N�,Ln_ ��Z�N��.��ѷ׏�0$���`�������?�T%��#�7�<��y|�L#qT	�J�~���P�X��rd�՟,��^� �u�}�$Gl3,���޻HC��-���Mɾ�ϧ2��&-|G����C���ρp��?~�Qi8����r��Q���tLo����U�ȸs`�=aa�b�"yB���)��W[���F庺�	�57��g� ���ga@X��,)5 �ӏ9P���Q����r���h�}օ�Y5E��dd��U���ζ
G�o�-:�4qG"(E_RI;�<XY[�Xh&��j����"�Dnw([�L���_-@���[[� �4S��e&(��v��ɹ���K������L.F���=3}էw����?���M.8	�, y��"DOQ�2'oi��q2�ᬇ����^+��u���@�]���ː��v����~�������t��9@�>��lqY �d�׆#8���{I�0��u����v"0T�9��/Z�GW�xiQen���'q\���8�v}
H�*Xl���)!�YRV(?1����!���ٗ�*AFc��4�F����T�h�n�V:U�n���h�v��b<Ж3[]�-�Z��-��������ڢ�W��=Sq@�>��%�m����aj?G|sB^����|���vއvn�Z�B��kc=���ܯ�����$�B��U��`���\�q!-�?�z�\��0�RZm�Ox��&�4VKY�aIX�}�ڠp���S\ԭ)��*@������&a��t�2��z�pEo�v��IJT�@�^t���<ҳϛI#`@��)W�x"N�Oi��T��i�qtV��t�A�i��,^^�U��J^�^y��ږN���'+�@�fϸa��IV����m��g.�h,R�ݥ#!h����� q�scuU��B��w&�r}$Bާ�]�2ZyL���U� � ]��3�^oP" ]q6?7��_PM���2�Y�sB&f|�f�� 0�����8��b��~9�Yb� n���w ��I�}�>�&��.�B�l���y��/�tG�Z�˕�9"N7�H���iL���٬~ᩳ��
^�$Z���w@p��1�(��e���+���NgY�B�WZ9��N*<0w�8�D��X���,Uˮ<���#���Q��X��;˔4'5U/���v(��Ư��Q5	O��C�a�Ԋ�e+�~�C��k�-��z��A�oH�,C^ �$R�u�]]V��+&S�"đ�q��o�� �\�s�",V��u�!��r>���a�v�����D�c&��g��y!�f�������L��z��1�mR,�]b�k�U;ң����q�9��]ԯ��7� J��얁B ��d�c^g��ۡ�Ic0)c�Q�Kn@�ɑ�-'��8�o�#>#̆�$;��ۭJ�-K䎑%Uc��+ض	���(���[����Z��*w���0A3�8�E�������抚�F|XwSI=��p߬��uX]^q�H5��\l\O���L傕��������[����N� ÄK:d�mƀ��BW�@+�Ƅ�qx��Q�/|{�y����o�RR�4��]�z$^Gus�|���j��Ed�c�@z��d
I����%�-��hE/���}���cN[X�3�������)DH)R�GIT�Ƥd���/p:x�C+��%�t�Q`Z��*6E�S��z��O��Y�հ���f�v���O�e�H�aY��տBQW�t�݌Yh��E��_f�a,A�ւ��7$���9�T]6��;>�{����S|�H[,$AϷ�r1��^�E��^�33|�p}�W_��Y���T�f��PO�{���
O��j;թ'�L#̨�` ���SON���oXP���ٞ�(X<�iI��ڠ�lL�w��K[ɜ�meY�G����pf^�r<�U՞+�Wү0>����o5��A��*�����O}V6���H��7?��.�GZ�	]��I <à77�sj�	����A�WJl�ԢO"e=��El��*�] 'K �$ǫQ��]ڨ�`��u�MKɘ���m�˸�k�(e7de�Q��-	/���#�%�|���eb�K���X	��J㫝��,�� [9�'k,
f_ir^D��N�n18���
��PAV>��U�����c@��d�!+�C�ɑԍ0|�[�+�i�R��ք{}�?A���N�m�Pݤ('�m����9������x��a����Gc�˲�p�KI�_{�S��&&�P�C��5Ɵ���� ��\��q�@�09_��>�.��)��:�_+�DG���).�s���|Iڞ��6��.�FKo��w2�����W�3�"�;i�kEK���8I�J.Ƀ]�'A}��r�r��d���]��D�_�Ib��Pl\p���L�.6�r����hrIjo�LPi�W��6���Z��cz�ܺJ*=���I6�4�t����V_بfé]�|+�i�er.G�۔
t�0)Z3�� � ��f/�{X���}�u-n ā�yI�e(m ������U�"(kqڧ��G��CkfLIjh���_�H>��Yֻ_�B�2�k!�m^��'��v[Y���O���O��εҙ^4�;$�|�\h���N���>��[-��h������h��{���Y:x)g=MM8��`�/	��#'ьO�����4���u����-D���0�$i�<3R)��bAxݬp��o����V��M�Z���L���	��.0�=� <�N��
]���^1|�qHN��e:yX3%M��cnD5Yb�	��]\Yلx�|���-�Od]����[�쉔�	Ǆ�i�������2��!s�P�k9�6O"`��q��y�J�$9C��ucͤmƅ<�h��('�&p�mi5����r7Pt��$�0S��&M��J�=��X���Z°m_����NcX!v�@}��"E13df���Kw�8�RDUi�փ�����L��F���$ȣ��ZΎ��V�:�H��T�����cƓ����P�B��%0��{��:� ���"��nF�+s��K˯��o>7;�d��c���6�ӸA�i�xT6�Yp�����Z�e�K���7���v�O*KU£���Λ�F���l,��N}����g����pS	�U�P'd�[ �g7&�,p`)U2��I�ɓ�"���� )��x����@�]�[�_t�џ;%'ղ1���l'T	�1��`[�Zo��0�#���Ϣs�����9��U��S��q��lN<� ��WV���t���>R��ؒ0)Z���g8���!ƅm1h�)he�~�a���|9����udT�}Ҽظ��{��
����I0q #Kt�K�������讦|�_��$g�=uy��LF��8b�2���t�j���O��GtE�j�Z�r@�!��p�R�Q3%���S�|_�0ޒZ�N�jڤ3/Y�|@;�M�@��T��P�7whP|c�S��_�����m�EKTn`��Yr�HX�';�S�����JX��d�M��fn��`h�Y-��z��S���5E�~՗��;����%��j�~fMeP���6�e�lք�t:[�P�y�9}-ŰB��T�u�R��"��_�SqC��	�m!#'���}�7��30��A��!��z�����C:�ɀ��>]���p'�f�"����E�J������4f)YW'��,�"��o8#LNuPB�t1-,�j����z����m|�."��G�&4S�a�B*�uME���g��/�D�=�1�A;����L�����BL�Ug� c�n��� �\�٣�~*Iy���Äz�*�xbcg�ղ�3��w:�BD�3-�rm�y�6`�T��3����?^���5*��f��ۻ�sk�G�V0u$��7\�Ct��G���Ʃ��ʇ׾��"��cw 
l���g��?�ެ�q�ڽN�>��Q	���~�\��a�	�Zw�m��S1���@��U�j�����Ĝ�êߖF˔{5C� ��r��%�y�Ґ5��fpu�>���)�q�-zO	Ԁ<p��LD�x{I�z���2�u|�$]�h�&�����o��r∫`�&��|�&�9ӷQ �ȍK׆粧*B]�]���$:k=KBʛ���݋��D��8��=<�Dp#��UJ�pe�<�9mfPo��1�n1I���m��Jͩ/�y���>��&��$I�h4����vJ؞m��-k�I� �Zya���ce��g�g��Y'�·N����HY��4��U�� �ͫ��ʁ���'��Պ�������.3n�W@� @K'�NY/�TR�����Ғ��T�R��)��R�����*��/C�%
`�˪u4f��5��8�X�����;A�wR���kg+
�;m���\pF.�Na'����b���<W���U�^���C:�*����z��t��1��(7f��^:�V��H�j�<���q��s�HLf!@��t�+r��$���y-�^χ+n�����XQͳ!�+��b�5a^V5c��LR(��bu�.��(אm�YHsE&��*�����Yh�f��oR��-���A��55��aHMr�ʷu\�ZV[��/8�2̳0�U\�:�,���ղ=Έ~i��ql89d�l�g76E��"�v����)�4����<�� �.��!��׹���`��滄�[N@�I~�:<Pe�{��n�(~�m�%�(]�B���~z,�#�V:Rg�D ����OF������_�I9�i�^�]��K�ϕ���d�k2���}�jBf�U��?(�X��8�{2BK�GǺ�F�R����O�I���DCx�+m�^������|!�f���{���TRz���[��Xg-j��;u�Z+�v:����F޷٠��F�Y�l'q��>�ܳn:��{�s�)���<k�(I�B�.�����#x̭iq����X��5d(I����E�8���+���}w[P��<�Y[|D������o�Լ��Z��2�	)v-�����z/U}�a�4�[Wֹ���Z�[�m��cr'�'�	Pkp��#�c���P܏}����/KC �� C��SՁ[V
��c�c�:%p���e��\��{N�����r�O	a���9���\��ٞg �suIa���8������/������ӑ��oY�	q����o����܀����k����M�ń/��v?y���w+1�C:B_{;���%��:�뎽�>m+���5$���x�=p�|�?,/��[0��q�
�����C3R-��q�<�+�1�0������q,�I&�X�!~X��-'zt�7 ���_�n0�ǡt[Ru(E%Ӝ&��E���D��.B3��W^X�<����H��'�F}�3�-9^_�
.����`�T~��$�T���Y��X>,[�=�}���iAw/��&ny(��l�#������/��i<�J��K�dEC�n��sUd<}��{T���w�Cs�(����7a%=��,�̺��wdٱ�Js����ڻ�`?u��H� s8ݦ�b��4��;!9Q����j?���Q���@�3X͗W��+_t|8�\���?i7'��Ż�6BG�:O�)p�����?�I $K�E��������8�h̘*<�����t"c��,XaFj觡'8T��]?M ��MW��6�R�j;��X�F96�)X�v<���exT�K�w�`S<4�q(n�ʮ�Й\� �#d|]��y���b]J�5����������I닇��{K��!�3k����ྐ���B��0V�| X�ԲZI$��N(�t�gF	d���7f��VV?���A�Ъ��@a�.�$���0��&@b��/�Pt��=�DOIѴ)V�uA@3�]K"��2���U/�M�<a�k	��F��p�����˷���=w�ڥK�������ü����4���E30�B�v��k]��<�Gܕʞ�T0�;��?-h��A���fI�"W��Q{	q@@S�A��j��~�q��Os�%Ȫ��� �iQ��� �����B�uf��3z�h �<�c���Q�Sb8`���+��vE�+���7ɯcZ�>X`�u@�
,���%��r���kC"M����3b�,֌��2����l�g���m5�i}��ҧ��i��m�n�C��� ��'�}�k#p!3 2�ȑ��t�I5�{�;�&��֞T�9��*����oi�\�
�I����J�B�_v'���3F�ɲ��<zI�֫~|3X�s/��/婈��	ZR����glXk�ʀ���H��;���"(�������/ك_��"w�$|Gl�����,zZ��b�U�|5G��|b��/+�h`Է��yY9x���p.I7Dt8ZCJQ�w2@6t����H ���0,�_.����"h;�i�4KsP�O�*5Y^@4q�qfh +��Ig��+����#=x o?�2�4�L~�f"K�"���IC�0�7r�b��ʄzQ�g�=�&#=l�b��cp���Tݔ�QG��]�zL��n�2,��'QW!i��d㿟Ԙ�<k/[k��v�+��za�NV��ߌ~��2P:�*�e��X�Qn,�
K�4�"Wf
|�a�z�n�˝�1U�^�E[ۇ��{�c)��O?(�jf�?wi���iB}��.C�6��q�r>�\ k�Kc̅`>K�}ש[�C�������Y�x�ȸ�Gk����&�P�)sh�܍�7�t��X��:��V�P?�V����
>Yjr�S�R"���J\���1~zr��G���Fu��G� 2��ɉң���q�B��
+N���Y]3A,�@���f/ì;�ww��Zki&0E���c׫IC�-E�}K��_�^�%��%������'NR��8GR�V�7����l�ܠM��Z^�8�`Է��9gv���G����]�o�4MiY���ÆL� >iE"�s2aX.��X��)4N:�7#�����/_��~m��^�����7�;3�'çR��X.�w��~�b]�ӗCU՝aK��Mu�{s /�R�m�&�����`� �E����g�n̺�큔/�Z����X�\�*�l�]�-?�K��ι��9������(��Y� &)h{(����.K�L�Sz�8�h�8��a��<��췝��z�Ҁ��Eb����0�|���v������zVJF�]WQ1mm���s�QFʹ�q��ޚ�+��_��r����n��əD�x���/��b֞X�u���ŷ�e��oa�0Tꈺ5Z'��͒.��<{$�</�����?B������vڂ����Ĝ��m�Ӧx3���跔؊)����_��%��M�������
�a?���=��l���r}�}ԘWo��X�(`��r��`�5C�J���m{����3w�\���y�?��8Ұr�,�H�X��T�!�� �*k��vI�V\�0u��P�D15���'�!x�y5(H��)�~�8�K꯫9���rvr�)�EaarIs�%)��E@��\51�i�����'5c�^Q�3�d-�Ү���>m�����ɧ����Qa����)4}����� ��W�"��9_
����h��ȭ�9Z�@��"lf�q=z��{�mݦ�	^��������(@EY7��^-�H6a:�f�����s��ݩ�v:{|�;��]lq�W���ٕ��K�Q0�ub���!��ֿ�0J�]�1��T�1�cPO�ACT�h�e�ϙ.�D��%ᓤ-��9R+8\��UzI�[�kV�|��� ���}̚�������A�3�H����3�[��7]:$t�Ӂ���~�W�@���i�B����B�M����Ĭ9������A�� ˉ/"��	_���r�tc�g��|�����~!�����䥈�\,���'�ٝ�'�Z@�כ�L�.
�g8�>A�{>��<�'�t�S���;��"�����h�O�%˰1��@C|�����`�h�L�Q*E̟���{� �ͮ�hbI{�]H�jb�I�7E�����ԀAz`��6��Iϴ�U���aB�sfW4b�y����\�����%��}֯��$�i�%9���<����3�f$��\��P�#�s����u�=�q����i[u]A�[��g�ȴ�>�<�k��T��3w���ed��Z�]��K�������M�q#����֝Si�P�j�ZΛ�5�T��`�c<���^\��
�%��МZS��l�%�)���%ֹ��$�H���7�b:�������7��p8��%C�]�O���ӛ�`�叐�V��ą�����"ٖ�fb,�lQoK��3l�-?8N4�7뛖���R��1��q�a؊0�>��2��m�)��հu�"	;���z�7�=�M�K!s�D\H�az����N�tL��b��W����V��ᆕm�[Mp),���_$���9�X�����WM�@s�	��k;�Y���l�+
AL�W����p�¢���5P�{v�z ����-^eb[eLp�R򞩩�7UG@�Z_��#�����|��.\B�h���p=]�\����lk�K���X�s4��أ3/�K�v��-_T.�޺��F��d������ٙ��뚡�<!����$���,/|�~�8Հ+e����*(��d���6��J�BV�'�SW�Yrl���h�a#��>zf2ࢊ�1z�w@&;���x��M)��T!��$,l�ebN֏����h�I��+�>�%�T`%�	(������I�u��)f	Z���b:b["P����|1IО�"qi���&��q/���S�����Hs�("K�vH	4���@=��ژ �gB�[}gy�pz�Qԧ�Ȣx�Č��	�H������hA�;�ڊ��9a^�t�ՙ35.5�f�QFtw������6�L5����h<"�.(v?<\	'��!!�
c�A�5����OSF�W "��N3�,;�c24�� ��)��aÊ�[:{Ol�m~sF��r�4ǐ0��`&[����FFp�iŭ�	'�]ajK�Zw_H�Ck���`��=0~�UޅC����!tpW5Ò縐5 �~�APX��q�Q�ԎZ�`E��Y��v�>�B�n9�f�
�U%�.[�c��˘��H*BQi���7�B2��ͤ����lWl{.k��3' �Ԡ�m�;P̭��F4	�B��e�ӻcou�}�[W a��X�[>�5&y�3q��P��:>1�;�V�Ftp�i�rl�!����/���-�~�&j���Ax�րQ���ݪ`���
��J�\G~�b<�)��c!t/b�D�J�T�Fއ�{R^�,��,�'#�)Y̥'�rA�O�{9��,��by������zx�6.6��.S�j�}I��pP!�lN܈㐋�o=)U3qc�m�r)OHx �I��<��o{�R9��FWOPN J8�y�����5]�B�u��ن���һPl�!g�&S�z~�
�PN���ϑ�:t����3�xR[�*Y�)T����_!oY��a,�~N˼�����k$ے��8N�c߽ǯHR%[��*�Ayʺo��tR:J����{t��#����l���&2S�}329)��p	�9� ���U�tn 7m_���l񕠰�<R��������u�,!|�����ñ�,�����e%S����}�2z���<u.���}�ۦ ރ�,qDA
�#��-��黋u��|�:��r+|]���ȷm5���`N :�﯂�~`lAh�H5��W�^Z+�
��P�_{[��RCb��l��lP'(�i�/V[[o/��F���e �\��:��yI<�~=ؽ���&	�a�9z7}x���n���X=˪]�n���O]��)W��4�w�K�ދ���s�O�;���oԺ��Nr����=j�����\D���m�*�9�V���vhb����N{k�m�g��CɄ,紙����2�g�1��[�d����b{��䩽YUeKV 5�N?P�Ł�忿q�ws09)aUM,=��.��"��0�n�U�5�P��#�����Pu���/~;�M%3�1�����܌/?E������?���9��n��z�+X�1`'��dBz�a�����n��S����c3��_r�.������D��RB��������E=�[��ʒﰄ֢��ZP�5r�i��G�L�}*�-.�ٱ~�~�Ƿ)2)��Gq��������@�a꜐�ex�f0v%t�+Q��W�F9�� "F��:�JA�����>��ɮ�JǓ�N�j��H�t��A,���U{���jƷ2^�R��1��Yp�Z�*�P} ����U�i;���Pf[�g:�5�`���B�	n���en���os��°��u���΄����!���B	Y"��8?���~�N���g�2�5�#���H0�u�`k�(���aAʖQŻX&�iµ	��>4��>,�{>�����;3Bc�~@���� �k�2P�GҞ>{���Ϸ����a�`�"�={B��3޸z֙�e��Fv��TΆ��"9�\ 7U[#��}��!��Dk�dM��돸�>�8�!�Q���i�9�O7aW�4�bS&@�f�	��$�Y��6���2`qo�c��+&��8�]�JEh����6m[�e���3{�8T�UMmp����M�3��6h�G�<�=�*���!"Y3���!�5۫K��̀��7g:��{4j���o$��C���g@�_lGNj���b�l���ől�=�pm���w��
,t<Vq[{d�b�%z"���KT0�<u����7�I']ɚ�ˮ���5"d�P~⬂%������ߦ�-0�)6_V�%Oj~�VrN-<� ��~}Hy��a���q�j�Ψ�NE3���!K/01��y5?��c|��QH�hR\���#�r�D���5������\J���f΢�������"w���e��ymZ���D��Nk(��C�	V�p1��غ���S:��h*4Y{:��^�$����7 ��NF�u��4�Y.�<?�"e;�KZ�G��G}@N�mO3$
It�#{���V���zm��C�,�����7���u~7-�4)~�!���X��9�~��-�SV]< xo�	şΚuR�2M�'f+?Dc*����\�kt|��J̠��؎"���� b|t̆F��C�s�fg,?��q����L䮠��@�\W����X�PhT�>�BCȑm�>�mh�Y��Ry�xc�%Գ���
�0�H�`�T���G��ö�]���^�`j�{��D�݂�����FkʟM[/�D�<��w������ ���Y����L�]V4X�X�^Y�1�O��V��'^�� ��e�q����?����=��p�P��Ϸ#NÖֿ�+1������@K�����V(�DBɘ7�S?aK$��W1��S��U5p��3�G��;d[��K���1<��7���n�;.`�wC���՜߷?``��{U��B�WW�������H�U3|�\Ծ�8� �h+|}�΀�ō��@��#k/A(�&�*I�7}��I�r�3��<A���IS�sm\�:�݆�����ZW�g�k6�mF�&��/��g�$������/���a1�#0�a�yb������@,k�|Qh,�5�;����V��w6x�/DIm߼'m?��+i^�0�2GJ$�, ��"��g�1�-N�����}�`r�����qS�R�LB(e�"B�{�v7t��e��-ݙ��9w�f�G����8#Wz�+M���8F�$LXs	yL�P<<�w��o�!s"�O��~�Q�F���/�,����D5Lf����f�DeѝEӲ�9�ܜ�g�������J���J���y{���m�HA�K7�(�z�/3�X����%OscM:���Y�S����À�|z3��Z6�9���~r��E?A%D�R�*�Ǹ�)�.��",uR�*���ߠȱ���L�w�	Jt]f��6�<
�Y����>D��`��Yn���a5k�N�:ݍu �<6uEŮ�&d�xQ�貽P섖��L�$��p*%,��ڈEEFM8&lngL̿�;����7����nL��!�&��;~�B�ʙ\���Z�_%$Wޮ��_��/V�@����e��H#��<z������isN�Ip���,��"��B����~&�=�ڑ���qRY��!��}�m��s�!���Ѡ<��Vu>��,9�TI�iڮ�� �t�P��G�ܛ�q���L� �{v����1L���[�7��Į.R�����
�,Ǣ�8���eQ+=�E§�
b?38�7{ȣ�U���8��w��>5#,{�F�%bt-��\ܛ�[���X7ޑD�]�m,o������h���S����y3�DeV2G�E�E,n^�˶�?���5(��k��"y�̓��޿��z�ӻ���Z�u��J��<��A7יּU���4�Q�,�TY���u�M�j+Sۙ��e��d�Onu����4�+WȌ�2G�a|��ªAJ�i��莧�'�Y]#Ct��q=���b.��}B!p0t���Oz\>r~H��$y̹z�O���_�9L?�+T�6�I>��Ǉ�3U#y���B�'8}�G��D}�v����H
w ��� �����p
 ��T��`Y]��<��'�Ջ�؉!����D�Ǩ�� [ęs���?�/�,fs ��zh��99��Ԣ�f(I�)��2�R����8%(0{�L��A���P/�K���ͪ4��נ����[�ҪԨT^�/��|������_A ���3���4N��n�
y9B4b�z׿�Ú^���S�ͷRP�L�I��_���v��^|+�_��ѭZ|Rpk�"S�#�>b�'�?sB�`q���N�ejX����N�-�<��;�_��}d<�)����e�C)�Pĉ|�Z��o�mmKeˤ׾�D/���/C�18�M�Bڷz��U^�=��+���F��r��� ��-�R���U�͸�-8'���c7�R������ ��Y�K��/Ć���@���"'�!�.��i\�PFU�_�3Ҳ��
cgZ�y�.r���FƏ 2�)ziq��2y}�:̘�&iU����F�.�_�ӛ���܄���oG됟��+������V��rշ�3:G^$3���#u,?���P�B��E�HÕUT��q�̍{:O�I�J�khH���s�]»-~��VL#�o�F=ɢ���SF�W9lV_�������n�:��[4WX�`�}\�ǃ�Ae�o���fV��>-�HZ�l�øl����b�B�A`�����<�%�)�MK�7����Z�:�r\Q�O�f�ە�)��h�D�势�}*�ΨoA�@=�� �䐓�GIrݞz}�(_��M��#K44a[�2�%�g��d��<#Ϗe�f�7]��`�=���&�:�ϱP�5��9��7�����p�"}�L�z�J˔Ш����z�m�.֧B���T�Eֹ�L�F��=�a^J43�^���8��j3�Qo����_�mr��34�䉇�G$�N<�~�$*��7*�涠�P�\t_��w�pɑ�D����K�d�����<�c�JS�o�
�X�49d�(m��oʷt�Ğ�f����k�G�2�"4��`�ǜ�����%E~�Y��F�*����d���ߞj��awrf�*��'�ðef����(�Z��Aٟ�kA���91B�2�	�7\�F�(�`��7[��o����8�� ��z�NUi���B���S���E?#��<d����|p6�~*��_��2j��{t�I��ѳ��z=$�twC?����E����Ǘ:m�ZY���v?�[ϵ�%{#%��:��*5��j9��ۋY�,t_�i�!��wl/q�vB5����ȳ9�ta��T��UVq�2!ʽR�:Ij�}㠟�H𳃣�#)�H[�ݜ0�s��	5o���2EA_��)-�n����o�+5����ȖG��M�҉4Z��4�IV%�o�G��,�L�D�� %K�.:�Ag$�*Ǎ#��p�/���7�����&� �sz#�5��g�-�"���W ~a����+GB<����7�ד�[��1_%d�ߕW�Q����D��kM�����m�oJ��h;Ue4�Eg*�lm��\B��Z<��V0C#,y5��,Aw2f����t�O oҝ!�w!�+�=�(�N�:�힇d��è�	��0��~�-�|=�+�j�KmN��-�,O(t�T��v(��v�A)����ɶ.�����6z�ϛ�E��`v�T�{��-~^f�A%�f@�X��������1Oi�'��xX�l52��CT� ����#RC�]�[��i���E�h��7R���O=��ڔO��`�\�&�%C_9��U��N��y
�|3�^�S��*A���0x����dL�?��A�np������Y�e�U1�	�cԶ0�*�C�=?oI��-e��u)+2㬖W2!b1�H��c+��+<��&�As���tF�}Sy</�J��a/�$꾨>Q��}��}ί�s���d�|Qy����s׾�;��;?�񯇯�m�gm�/��Z���>LK�ѵ�J��?Q�t%3C�fJ��lKP�C���ك�!i�|�KO 
Xr��㬲t����Y�hO�Փ��9�؝��f���D�B���q��8��� ҹ��%�$)�y�#:!�e�XG�I������I�x%��0� ��~)������z��H��25�|w�/AԬg���F���p����! �%�wo��o�z�0J�I�ْ쭸��zj�o"S�j����@>�wJ*A�?�� ����1v�.3��i��k�Q���m��I�%xz?�O��.��t����M�>6���Sr�a	���Mï��Ƌ�h��0�K��B�7Eҩ4�fJ�|�de/��� �e{v�#ɴ,��E�y?�9��ռh���%y��K�V3���1J��s�s��P+������c�Luտ�P���!U~*��ar3	�6�Y�cRLXl�E,��� ����z��� ~�C'�w���}��O��n�-���(���ZSzYN΁�o�e8y�X�>�媔��*����p�-�N8'�M�Pd<��l��g�a�l��N`�6̓��X%�uNd1
 ��C@��
ʞd����)�f�DF�D2贻YHQ����w.�ฏ���%�0��vj�s�Z���Zoi4t��1��2��������oF	���.�iw�Rd�L���Ob���Zɪ[^:�f����(;����*9Y�u��QQ�B���R�a���[%~5{�i��\��֪�G����*#^�=����4�gO�C%�H·�.�ӿqK)H�_�[M
>�Fu����d(���#d��~�мU����'^�Lx�&6�l˴�hf�{�g7�'�Uf{(0-�܍t@А:.�QcC*DnI�Gfm�e��Ej��df��W��3�����9��v���N�^�x+��N��T�5lky��;�|�|�Kx&��~���l{ Uu�>�p�pوIٱL�&t�3>���:N���^A��ܩ;�r]��W���Vj|+y��ׯZF�=�mQ"�ׂ��~^��4cH.�׃4̄u��WB��&�B��?�����8ׅ_��3l���e��t�t��GN9��bX3+I�#����%���ă}{�P�����mk*���d��K �ʉ��5z���/��G|_B�:�}{��߬��H~��F�uo ����K(���?-���Ȇ�ݭ�y���s_V?;¸a��vd�3���Q����ei����W\sGҧ���|]���x�jM���!zm�,d��su�I�,�Њ�B����z(K��VVA�ǝͥ�-ވ��zuh�lP�cO-,���ώ��1J|k��6m��v/�K�W�V^:Rp����D;�l8�TG46)���¨��~S���TE��
��a�_�����K{ۘ�V�檢Cqq~Q���7���^�iJ��C� u�ZSy.l�3�����}��a��J"�|G�=Gҋ��������}��G��y�� p�B�F��Yi����O���B��0O��5�q�l-G�8��-&�����e,�pu4n�AS��h7�B5C~H���� ��S!g���R���f���bf�@���v�mҹ�_ߤ������ߊ�sI�����p>W���Ck_)�#w ��N׌�V[���i焭������ٱ��)�*6������+f�M�lHy�/��nh����.���54�m�Tv|�1���%����%%�L�,惦�l�n�$�b�"%�a��¤�ۥ^����ܡ��tƢ��%�qLl��`�h�;E?�kAL��+I��uzά=������BH{6�q8�l�2�jVi�)ޡ�
�Q�`*�i�!-<���A>~���\]]��NJ��_���ѩ�n����,�E��F�yU�'�_�_s`�t!�`l��m��W�����t��L��bQ
P��	'���C�z6Mq�j�iY6`�N8�5p��\��>�G�4�� p�[�:}M�N�ı)�e�T6��U�ߔ��7ޏK�>���B�*��z���(Q%9=�rz����P�hJ\�OE��ѶX��DKk���<��KGD<�=rP�V���Q  ��JK��6n!g���a��'Y���T��㕟si���|�q7�����#��7���0�2����$��j�9�j��6�;'��'��?�J���>3�w��E�][bk�}�s��;;�.�Xm�j��"�B��n� �Z����:a{�6�Ճ8_� ��������X5e�>F��{	���ۚݶ)�h�Pl��=��g����r�-���k�0m��z�Y-
�����0���xx@�q��ٌ~?�D+�A]��R'�E��<�f1 ;����Ӊ?���J�;J����_1�e���~6����d����t>�!wM���W�7�7 �y�C�면��sv"�G��v�M�C�YFq�8}�L��n���Jj�qQV�8���G�|b��k�Pxյ�)�MTM�N����aԦ�ɒ���_�1�̡L�[3i��|��2�R�������C����+��α��	1�2�Q��Hf3
@�ɉd
qk�T�Z� �*�
qX�m���6}s���ʵV�G �̉͞I.�g@t���k�����F���9y����`a����a�Fxk�@Id�3�"�t�H5� VӰK[��;d���'�h:�S� �A�F��6TK݂<����}
�2"JC���X�N� ���}P�����?�;¸�OuWZt��E�&l0V�*&Z�⥴BJ(���q#&Sٰ�^����?����Z[��	8��R�$Y����ƘZ�a�8�b���/V�@���9a�L&?[O���g��pT���9m+U�(*`x�˶M�6:�7�[^�m�	��nLE9����lG�.�ǹs��)"����
����D-�b���� �8��e�bWǦ4_�ӡ�a��_=�8}%h�ƹaO]1�Z[�Ү_�����b�4o�Jm�߳��q��v����-0���j�?�[H�I��$&��K���
�� h���s ���Op���\��c���cn/�R<{����
7��ֳP$c��j��u��-�9�@)<M��!l�)��\�рq-$�9'p����YIC��v�"_�����;�5e!�pCDϗ�3w���)�y���������#K���3�X�D1��;����c���1&!'�I�(4�J�X�9�F�z�s<x|�J����a�qJ��- [�T�{V�&2j�0�5�4�;1)�J��߽�T����^��2c�R�O��q'{[���ݳh�a�(y��pBE�"Yt����E����a�<n�*夅"�_咥��+��}��I0����4�̜;
'�i�J����N'�ڑ��5g�F�c�6%����-�Թ�����g��:��B�������
�ғn{���F7������!�dݭ�~C۶�(DzgP��-����#C��Jïہ���#cFfV���GS��ȗ<q�װS�<{��4[&:��B���k�w~�'1���g9�V��P�71J
��אV�~��4}��{�W3m���H�K���3A���^!�b'F(�D��y�v0�=VVJ망lQcu\j�m���4A��K/f���sh��9��m%]i'>4@e���1!r�oVl�
r�`�ͼ4W��O���V% ��/�Q[Q�eU	B^!�=��|��Ek��	�{Z��N�,Zض���2{����u�h ��5��"��#x�����f:q��]ߥJ�ʇ��6n����I8�Mr��di��@�#�Q3�"��`���I�k~Z���;�7�ɂi��;h�?3-jT�t���B���Ai�VLN�J�R��ʬʟ��������nEG�A<�C�h���ő��D}��f� �����"�t�qcG�c��U��P|.�Wl����w�梗���=:#v .kP>�4c<�v��'�ߣ��Ev9g��h�s-l-u�k+��L�ޮl�_]���xe���q�� ��Ś�_Z������in%�k�098��8,1�e9 ��:�%W:��,AsQ�،��g/^+��o</��Ūx��@Kd4�cn$�"uI���k
{��i@�	R��E~�[v�)�n���=��}s������-�Ux�d�M���)?��[�왣����*�
<�4N5��O���Qq
.	U+Q���w@p�~p������t�kP�/��&�iF��sǊ}x�qZT�{�od� �"�{�Hm�;|,tQR�oI�������^)p.&���D]��t ބ��v�����%0D�~�J�B ����j=ɞ}��Hv�j�`������t�-XAw���� ��=���&�L�q�y��i�A��m�Ă��O4ϵR��
��(�:9�ܙ,PVCu��A
�S�XJMѹ�3W���|��9"Tu�L�'�9�)��eU&��a���y�����rU��hȹ���ψ�3>�	?P����fH1;P;_4H�FV���͙��18$�w�X+U|v=�e��a�a�4�;�_�ݺ��t��7z،� G'-��mXx����[7Y+�����z��&����$HFa�a�@�mB}�p:O�5?���P[*R�IV��dL���� �B���~�#��⺒��Cu�>�;�
�H��9����#��D!^��e���A�.+Ka��ˑpA�BG��u�G���ˑN)��n���;zc#��δ�f�R��	�)(���v��d�[���$�x˭�V�u@�G~"����8�P"�F�yRg.j��ݢ��0��:)���V���D����m��V�iݢ%C�p�6_�*��,�髖)�������b_ i��%\�Y�# A�39�R'��b�T���Xlm��TE�ɺ5\9�/[L7�o#�6rK��G��;k��� ��=Ey���ɴ½�����_��5����#}^�E�.F��f��'�P�Ғ`���"/�s:���7��z�
T���T� 
7�qN:vS$R����
����JQ�q�i�( �1w��
Pß�4lYk?���<͝��O�Lb�����Y��
1i�Spi
 c	g�@�f5_�{����Hd�����:D�0�t��:BW�<���i�]�Oy��R��f�,/�9IeH�V����#=q���ՓH����hA������"��ٵ���2|��N�^�xwz4w|��X2;}(0a�1~��'����H����5E����ʂQ��N������5�t�?�J�әG�'�T��h�9���0�}��3�:�Δ��	Z�ߨJ���5��~ňߙ��:�Dx��ـ8L/ͶgTT�`��!{B�1�*��KH�bY럢�Ql�U�=�g��_����^0��M�0xc��(�%�Kz�N�+�}�%; $J�2�d��*�`����iC<CWH��)����a8��/�Vh�v�3�q]�yw��sm�8�Eer�ƌ!Q.�J(Tْ�W4��n���]���6�]�{o��;�w�y�o4�PVv'����WKx9�",�~�x��ќ�����u���$��ܵ[��/�	W�c0�k����}�,F�qe�hSc ���.P���E���(���d[si����ƏNO|W��9�E3��H3�q8��Ή����|��H5�`;:X�q�A���I9?ʛ�z�w/���z�X,H����}�@���I��K���@
)ۂ��r��tTv ƴ�)R�!�;`u�]h��yb/�츈�{�˻N���ܹ���ϴcJ����I�T ����SX,k�&�?{���gl󉂦����M�����[:�ݘyy�5�ڑ[P�S���R�v�[Ǐ��@��Ƥ�L�h�N���\לu��ML6�K�=���]�kb�Eo� %�1<�A�i�y�Gb��� ���|�馣d�
���w�̒BI9�{�8���P�s��E�QK�(��_�/��q�;��HPuRR�oM>u�ܯ�蜂͢�����TcZoNX_��Q6M�҉$8h���=?3�
t% ���16&��,�Lҁ��`~�� �VQ���}:F]*jIc���m��u*"��t7P&�l:m�WB�+�d�I	����2�5��k��o���6��O��pX���SU��p�-*��c�V�Ņ�d.>,W�.D���ҥ��-<�@7,1��ѓ� ,��̼���f]6�/1�E3ZeoO�Ѹ�T���N��V
�f*�M�3�w��A�	�=[͸a�O�����1�b�(X��T�StmoW�h������#%�ڪSy@��^{1^by��f>�y*��l&��zz]�2kS?�"�*�LΖ�i��R�G�ր�U6i��<M\Ł>�h��"!y��g��^o����u��Z�\��l��Jޣ���r�=�b��~�R����Y�$���K	���à�J~̇q�!�Z{��A:�BP(�����D�����Ȑ�Ʈa���l�Tӳ	-xY��{�Zm�8`~�d�.�=�Oz�T�\��<���/@:����b��8�Z������>���r�����6RDz���z?ၾ�m0͢���t��I��ފDa{]��j(�wVj���,�>�s�g�i��>��aU㗥s��n���_�p��������#��aH���p���S[I�b2���,��hR0
,�x�EG���L��x�p�y��qk�Q�wL0�b�[��Bd�0��O�_h����	���3��JwF��H*��/Z�-�Ѣ��Z��w�}�E��uӆ'������J\4ʇȞ��N�(<��ȱ��0j	o�+�[$�����o~��gl$�QY[����	�(�
A[r]�\����*����!��Z"5yǂ�|�9`�a;�l�i��$�Gt+V��vE���r;Ӎ�K.O�bi=k	�p(�yq}���nr	[�����D�i����gj���!o����v��5��0S��˭$Y8��Qy�0H�Վ�/0�"G[�H{V�-9�Xy�C�o���Q����d�݆�#�͢�  �F̯�2����g���2��+@�2�"�Ă/n��"R��<xg$�`�.^%�z�\c��G��y*��	�8�E�a>4_VQ�`Gp���Z�@��_�+��Æ�*��n0�Y�$T�� ����4+�ƍ�S�:�vd�g�.��u��',�����%��~�~�2�K����&�j����������NW�N���<�~s��,�3�ВX_`��h��O��k"HA@A��z�C��T�%Lb�>h+���[B	Yp��'W��-��Z��6����VO
�ܠgI9荍 �1Ϲ���x���{�me}@����+�������$)�my�ޔdх
E��L�E��!�����&D~U�ߠ��o��{�_9�^�#��!�S��щr����+A�,������#	�+`R�x\�trd�oSI�/�AK�$�+p��[����j���_{��\_�5����O��A ������]-��ڹ�%GWKs�~�t	��N	x
���p���eU|g�#�8�2�a ��,{�w��3c���x�!_(|K� �Em9O�`�M���B��y*��r>��&�>��ʭ�L%Y7ݑ.�N��b��H�F��������lEB#J,��EX���[F��}��>7q/���]KK֕��������[p�u~r�l��q�E-#�22�B=��y�|�8fZ��������5R�t��eeQ��p��,e��uB!��10ބ�k$(��=�~Ì�̏XRK��k%���?����\����zWLM�T�Eb�%�NM�Li)C���Ҝg����vq�si"�)y��e�e��X�B�B���$5'��(ro}8	��Y0;�����W��R��g҄�/��t:ƍ���W�iF�N�I�kj��KK�e�dSz��BSA�2ÞIY����	n����3)��U��"ZC�~eW���㍊�X�L�7�!u9�V���{�V�ǝ��rldt;i�y�M�9��@���욹Ah�lQyM�����+��R����X�@~&1���.>l~�NՌ�z���@WX�L��#���w��|y��M��5�c)(����� �W6	^Mz^�Jp�D8���@O'M��V�Y�Qǯ������$'���V���=s��N�lJy`/�3r���DS�1� ��k&w�
t:+ɥP=T8�?ϗ�a<�@H��_ff��v���"������т��i�Tf����G��Y��;?7�� ��c=�h��3^��SPy��k�P�l����j��h&�L!tfI��jOۮQ�)YhIY�[�mkZ9���a6��"�>{�lg[�˙m��8���3�2M7wC����)��xhm��d[��>��R�l5X۽us�����ш漣t���MR&-��61D�]wj��?VC����UR#�?NXX^T�C+;"����)���	#�,5\u�V�?V����db��?��4G��͂�{��"�^��H�	���j�r�_)U6���FK�(���c�ԥ�Yڗ޶f�����X]r`�[A�l��PT���c��y�.���'s���JDT����q ����Eɩ<�	�D�7�?ԇ��o�>!Ó����|�
KP�;�`Z�:�Q�(�եέS���� ���꥟�1Y�O���1��_,7�|�b>6��'������A%"�M��*(�������g�s��	�u�d`���,��)�ם��S��{��8��p�Nz�><���7A]��K�
zߟ��u�=uJ��R[��T����۟�)�ߦ�'0�}Bp��~d���ƏBb3��n/�G�_���ץ3��cI��D����QT8fj?/hn��o�Ka�~�Z�Ҽ:W1̥��w�]YU C��~�<�[�nnǛA����)�&r��h���&7Y?�F%�+P���lP��//FX��*��Jڱ�?�9�p?%��=E��"%�t>@_��;�+���I��-�92�z�F�#�Մ��$���8UX��n��	C�5ė��yEH�y>�e���&���dP��r���4W�{#Z"A����6a����.G7�{����Y�#�V�&1��1l��<��2>Q�To�5.����<5b�C���Řbiz֥p%�GB�!�0���,�+m���%<�����r58�����ʄ�G�E��=j:7��Z71�qL*Qm0�wFc�̕v_��:�Loʏ����Q5��)�]B����:^�В�s!H/.k4�~�#?�c���st ���<|��-/�U�ѭ5�b����@-�A\�m���+cF5���E;�9I��4uX.5�ܗT�B3��@�ȯ9���;�rV�l�ET�O�������⻁&�'+<��)0�V�ͭ��P_���_]'v���+�ȃ�cL���� ˮoi,�5m�l;�BE �o�[�NM4!����~�b�YeZ�ͷ%�D��#�R��bxC :��A�:/��4^ 1���7�̓����	����Q���<?��sļJ3,Y0C�H@��	c��	�Z�6�ّ�E�<}(ZY�[������b�K�!)74��}�1D��+��π:g@&`�r}���=���S�UjAaFh�E~"l�q��:�R�Z��T�i|!���qogC�!;qw�p1�R��NTw�<�����յXŴ��c��nf!"���'�Pz-�Ag;�}-(�Of1j=�N%�����ӿ����B	I8�Z����1sk@�I.�11x����8�퍞o�2@J�?��4�8%]���S�&�ܴ�]x�������t4$u~���[����� �����F�>���`Ѣ�w0�"��/n̐�� OT/+|�s3��;H~WQD��	QZ��'.�.�����xKc��ӗ�Mּ=~A��R�|'y斜�+�V���������rk�Jś��3��"�$�2;<�H[6���g� ��k/�7� %>كj�䶽���?��$�r��`P��2�	�ܨ;�B�*cc���VZ��{�|�|`�@�$'�=�� �F��8!�3 �l���4ͭ�V��7�?���7�YR��\A	N�R���t���^v�DN�4�=��!$�[��ոk7~Q6#`%���p<��)��N
dk�R�;n{��)ċ�8�\8��O/uL���lw軥�C�����pL��a�2���@<>�b0:gx�c��&�G�A(�o�➰�Ǘ�V���Y������2�	C3rǂ놁)�χ[��9�pp{�\��퍬��?r�<�����fE,S�֨�:+��M�?��pd��[�)��@�fV���>�K`���x�ZNy�@kO휮ԃ���=�"��;�Q[3�%��yVV$k��� a��R	&p�qV<�&R�B[�V�;O*��*�����<�/�;�.���2�d�w�b"
���Q-��ڪ���:�u�w��:�^�-à
�RS*q�ܑ������=��B�j�# ����~= � Cj#�Ƞ�QV=��ٶ�Z���7莬���T���{?��:�����2��^��2�ޙ_ �G���,�2���T���"f�w�#3���k��J���J�AP	��K��ܻ�w���C$�u��	)��UD����'�^�6�� ���ܵ�^nߍ-�y�2�K#I���nt��ْ1(��?Z����?��nJFOjZď�)���*{���W��z�Fk� ��h�+��Ԛ�|�� @&���*�Ə���k�TI=S6dc7��ڲ�G��`�
�g�����X�)#�F��8�#����<��@�b�"�wF*A�9q2�&v5/����ǔ���z�RO�_F�
�v��N�� �-2g��+��|�����:�6�}oD�n��� ez(>�/���4D��K��D��eC]Q�eg���aP<8���3�������Y��z�W��I=�|�Wje��0�����G���T� ��ޭ��gc�o%�l"ޑZ�y�:�T��C\��M��@.���� ��ݰ�����k�`�>�p����Է��[���U���|�`	��u�hJ�լ�xj�c/�0)M��S#�Jx�oe���W�Ҫ	��
�	eѾ������Yӥ1�6��(c�͵�n:��}i�썵H��+���zf�6m/l,&\7����6���%h]#�Jڔ�#���o����B�U��\2����3�M�0>Y���979@�~	(h΢(WcZ�̥N��P�2���?>+}��Y����Y.���Q�T���j��]�;�&vu~�K(*��"�X8�h����축1Z�Sn�s\�d@��o*u��W�;#k�9&����0�s��)i�@K����3y�q�k�9�!�-��e^S����ؖw�ǚd�Ϭa�\N�	;���d0S�$�?�t�$���`twɽ+t�	�;#:�m4�Hb��q��M��Qu�f���
��8�m-w��ؔ^�Y2zo�L��>�f8��a���%`z�@��B�L�azW\$�֍�4ˮ��9�Sp�K�[�X���ɧ3�ct{�o<�����9�@Q��0B��h)��?��Ϛ�����Y0��-���sU%����6>r�ҏ��.�����T���un��u�:�ˑ��~�v��ڗg�n������%3�� �m�<L&T�[�Uw� �㟑�P���]*޹F!2�,��u/A�5Z�e]^`��KN����mզ� E�8�+��ײ����g�Ɛo:dɗ���`��)�a�%�mqc"��c�7���� %�s�8c3~����B���zC�p6�5o�4J�|��#|F�Ĉ��`zm�!�f��}��	׹�*zfÄG����u�W�k���+��$����~�.���#~D;��-�����)���x3�E���/�8q�>���@`OiR�K��ӝU�؃-�[�k_"1�0�X5�B���(�~b>�����/_VEӏ��9Q.l�J�N�����v"�F����'$hQf��rnvk���h{X�?Ga�����ߙ�XK�����z�8; �(�q*:%L��	���$�q��F�>����z�s�կ_:��//nVힳ̴��'�Am����H�ѿ�hr?�P��	�Ӿ�� �B.$���iJ�!�NNg�3>��@�ʘK!� Ң�r �R�zG��f��_t2a�Q$.�+m�7����
.�=Fθi����X(���q~ n�vˊG��v��p*V�>��Z��1��˗UY�﷉��3}Ow|i�L`t�`/g�z�i�s� ���E�xZN�|I�3���	Ic�^&������d�|�\μ�A�&c�6=�65`��Hv��xA=�>s���`�m�'�}:�U��<^h\Q��W 6x��g�))��ڨ5J��� �*�g�h�b���Q�"yp��v
	�V�za^����XH�r�������N�(�0?ת%�Δl��a�+@L��&�̪ ]�J�E�:<D+��ph�������+2x�د��< Y�>E�/.����ڈ;H	g��*^>tr�������� %�fM5�\���f2r�T�^����gH�^�q"E��[h����M�(���\ ���qn��W��kȥ��*�U�b�YDx�.�V�%<��y£E�`~�ˠZ����u_a�o��(/W��d�d�d<�5w#��P?5�흈�Mq�� ��M��I*q)u�@/_qJ
���Ґ2����*�)���L�4�2)�s�d^�NpPh賝ۡZ��k>kf�^�k��v�B¾��L��s#q�Ոb�2�\K� 6{�bOg��6Fpz�!�OV�ЧZx<˂@&<�E2��^"�Y�кC����Ѣ/.Z����O�:q���Uc��F@jR��>��q�c�~A�߀��,�<�GQI���K��q}��^����!�z<��l�~J�.�;>��X%2/X�f�e$Q�]FX�K��#Lz8A�.T�ίfe�6�9�_WE�S|�d�+s�,ؖ�^d__�M02���Ӫ �iXy2Լ��\Ş&=��,,�����{�\�u���'�cd-^	D�u�-A�o��ʹ���x"�+�sr�?_+5������}�d�=	�v�`�L'z�����ʶ�Ξ1�5F�l�y�`L�t�4G�E��s-tML+��,Ջ�@	"�n,��9=���%�r��Ha���Yf"r�̳ ����.i�6��T{uA|��X�Wo4\�k��2e֥�,�߃ɖ��L�]ɇ ���d���_PfFk��M�H��Z����q:�M�Q9�D��F\m��P	B�����e�_���h_	��ߜ߂я�]�l�y�mY_I�2���� BH���l�4�~K��V�=��G�ڙ˞۫"����q&��9%g0��$'��������~YQC���PCGs������϶���G����ta��@��	� ��xe�,���1V��'aJ'󃜁�O����v�D'D�����O�
 ͂���fշ���?�C&VIĞ�I���e�=
��6;�B�?_""jj),�[�a���>�şl�RN
����/�k5>݌�Q�S�V�G4�נ7>��lmc|#ee��K�	�L���g��ݐ�?��Db�D{�h�DW�h?�#�'����l�um���-B�Ɇk�Kn�3�P#K-�Rk7��f�yd ���m����!�z��A�����r�,�n�ϡҦwêi
�^�g�O�8Q��Tk��ނ���h���gS]nS�˖�y���8.��Mԭ^��(�zb{��|r���su �Z8��-�^��PŜ�$�Ȝ�֢��T#z�N��j�!�Dg^��Y��v�L��WH��.#��sbCo,�5A�n����v�,�� �����5MV���?�t�Pu-��:u9"R�v�s!��~yL-�-]�q�L�<�/\��*�����l��*J���?-�����M{%zo�M�{��+��X�8�|e��]��`X�1A�p��Ʃ*���^穧v_S���57�x�u�>��	O�2�0ޛ`\�2 �v�6������&�{ I����y�V��O
�ṵ���掮�If���0w��>��������ǤT�ҿ[v��/fdk��|�mF�J7X��l���Á�Q���
�����i��RX��S��B���H!oӾ��Xe�WS]�
E�Ģ�p�<�< ؾ�DAH ?��������oU��it�Q����/D0Y��N��?����*n���G��t"�@ ,�h�ͷ�
��C���ZA�.��y�R{�Q��N0B�N{E'���^1j���։�C���m����p�=G�⊀����	���!������'>�6�C	{�ni���M1<RgĖ�|����:����ڜKdw�G׌W�γ�/hKo�����sa@��mK;0T���QBw���I��@K7�ɭ�8a�.���f��MvR�.az@��M�X?�Sp�"��ZVí�V�`;L_ �R�H�܆�z&+F�����Q��G�-���s��'QWC�%��@NT)>�J��Q�ؚ&��Wm1�a\���B��1Oư"@Ҷ��3�8��>a�e�]��~����"`�]�yY���t��\2_�����Uk\s���g��O�fI)j�!v����I����^�..Z�H�D8�{��J�'p��P�}u��$~�A�'y�Q��ned�|�vzv�����]��lk��� µi^�T�3D�(��(PkHW4����81Z9"�'�.<�5��/p����g	J���$<?@�\d\!+���?�H���teT7])��8L�Hdd�.I�: !J������LX\>l�K-R��]/�w)�J��f �)��~�&;1#_D�B��%�A�Y �w4�!Q�K��췛u�a�����L)��行$��I1C�/J�`���~�i�Bʰ���B��b��}c��q����i$��ݟ�+4��1�·	FlP��/%�o3l��B��X���(d��k���XMV�ITW�evk��i���8�)p��[e��>��p.�K��%M�J��i���Γ�A*��ϕ�'t,�k\4m�������8GM]���%�U� ϯ6�}S���-���|�bY ������^�h����{d2Lz&⽔	�\'�jpS6*6[�W:uzO�^�����Qb���t�lgո��5A�7�x��;\A��f;!:MG�!�r4+������^2r��*󈦑���� H�+wY�c���eD����/'���&�����TT��\�9�b�XWbQ��!p���������T{���a[	�T������f��O����|�z��8!8$~���xm��^���Ÿ-b0����ȄI��/��Ɲ ���&�����D|�ɜFr�=�<gL���j^�n$=l�*����� ys�Y���iڗ������B�EN�癲tJ�,�Jf�@�hO64��)�/ػ��A���(����}�c���0�� �o��2��"�ܸO@Q��4�MS��p]>d�k�}�Q*V4D�A���I��ܒ�d՘Ӷ*�2��#�b�X�_���]v���ڴ~�CtX��p�������QI�o�~��S	���)�t�Ҟ`ߖը���.�>��t4��2/@em�����ʳ�τ�4��>Gi������@�\��m-�G9u�	�?/���	C�1H�%Gd-z[ 9%� �I~����>}2C\���sQ�бdF�b��|��>�k�=(��a�}�|�����"T��e��0��
�R?0���֦ع�'��U��	=���1<7�({-�p~x�H���(��78���>��X�5vH�#ڦ��++�F=�ى�B�����H7��=�6�OZ6�4*C�Qy3룞�ֆ3�p�H�wi��9��|�Rm��!�_R���>	Ɯ���v:�l��K��\+ t�����8�����%�̠`�Y��4���¿xIzk��^;�q��-����[�Ѓ?�9>C�(��tPw�������}��g�s�9cr����,��o3�nB��V��D�?�Ϳ���� h����A�$�m�Df��W��+��3�'<l7I�xS&9���"!�
D�X�R�	���|V<N��x5�L�O����V�����3��o3t���&�l5�k\6C���[]UDvp�Yܩf��Ƒ��?G�2��\1�?��E�bW��U�جj���V,�������9�9;�ޚ��X{�+���>��V��3���Jj����T�FƷȼ#�_�H|4t�_W���������gڄ��^�%���\��-�V��o���E��vS��vnUvru��܃I�x�O��`?�HO�fõ|v�[X���G�]�l��U�֩�gJ}�՘�k�v�U���<�w�-͢���#.�E����M3� �*ޤN�ĸ��Z�ё�U�+]R��r�G?ˁc
>���?��ݹ�]��NDK�p�`���6p);=`9����O�3Խ'i��h�rR��^7�S�F`{��jv�"65p㗧)��@��%�.3�>ǆj�S�W*�G�@�`� l�=Vf�2t\�pt�znW���Y ����ԛe6`yw�+�j�K�{Ԋ{�6�Y�uI�)�-��j��z;�xpq�����[)�wc6��M�>&����١��h�Ґ���3�_<��@:r���z@�8���Ҍrql�ͥl�H�/�D�����;��ǼK ׷�ޗ��2N�f˓�{:�.[�ײ2�BG�}�E�᫲�xJ?`�@s�6)���j�"	yEݿ���]K��.h����f�$
���;s�-q��r;uu���T��'qT�8N�6)�ڧH[�X�Ͻ��`�ʇ�`z��h�w�,�%\s>	@�JECrV���@����l�Lfs����]`�.Z@�jJ*�����~��(�Ū�ȎQ��|� �-A��k���5�y���&�0:Gr���Dw��Ҽ�?��߼v�B`��ܣ���X�Я��*�)Q��`E}f"g���O}?:Q�-�b(�;��Y��W%�{Kȯ��i$7�����+د<��_)�hK�����Wd����B2bW+��)f��W}�7�3��D���ќ&��.:�**dL�)�hHQ�|Y��+#�A'OS��g��$����9D��@)�ic˘��~M����-y�7o=y�>�����0�\�h��X�YN��"C*�{�Uw}��y�1��h�m��'���ܯc��S++v�kH��$�o����o�Z�.5m����4�0��~'�b��E�
4�Xђt�ERdg����o�Y�;��'8�
'ʢ�������<[KIfu"�[V����m��LJ�h@^��06ԉ��D��L�����8RY���u^�~a��
Mq�_$#�++9+y�S��L ��T0�Ɔac{��鹹��+
NkcXQ5@�>��N�H	+h����b�-�	���mKe��Q�~5�=���A"�^���,���`�v��&�r��ɠ����+#��c9�4��MD��,?�ĳ���nWL��3�$�T
��x@غ]M�����f���O�� O������E�0/2���j�-B�����r��;��@�|�C�ϴ��&̯���A8��r�4�x;�7\g�8�u��W9��&i?��t�uuj��z^���o�R����fŖ�6!�^����ŝk��!�LW\�o��(�\'�G2 z�v��;qDED�&���F���?O�$w�x1�S΁����6�蔾&QW3�u̽.�F�79�a���]��v���dTjr�¯k���u�J��ަ���j��7Zl�C�1�]�_�Qfmh����R��.='�Qw۸����o�u\
�ifHB�����v�M����������T3`�T<��>L,��D��d��#�G��b�ռ"���Bw�02��Ǟ���lД�JdExM���3ԀY�z�����)y� ��i����Ӿ�3��+����:�?.�%��c�F)j����kP*� eGV�!C!��67pj��!��.�l��bC0Z4�9�ec�ҡ�E1!+�V�&+�7�|���(��AO��#��o41H�p�o"��GW	pQNI���eK`�S&\��)M���~������B��(x+(V�#h��~TS���:,�噩}�t��j�He8���1�S���yF������A�6�#�o�/��=���n�J���%���#��m�������0� ��*����K{�v����m�� �����ʀaSb%W�kR)�����'l}|�-1���X���A��K/�"��ᢱ�b�K!|V`&�����N�����9�8L���k��?�e����Ε~������qB���IDp�ö�'\^����4�o��0fB������?3�[)A�4Ԇd���H���_v�_݋s��;�\�����xT6Yf:��M;�� Sb��+���"�b�JW-���a�ݭ&��54�x{;�6�
�t�[*�}������v�b�L�y��P@�(��z��8�� P�sʈak�]�r����`����{'������ϋW��_��Dٜ:�e��a�̛�\\�ĘjYG����h�r�*II�+��2�w�ѥ�j0Oq����(�A��G��G�B&4O%�?�ߜ1��ew��ǩ2�!�S^T�d�F
�C7�/��815C�,���p-�,�kb�������[S��2U��)�#{~�BK}*T/}Ϻ�6b�<�"N@-�¹+i�qr�%H�۱&��^S
E7LՕ���$"�B���J��UEfP���q�7vF\�qJ���}�W/�j�I�� >J#"i Q8�i��G���bFˮ��&R���C�z�<q:z)�.�Ŵ��Im�ќ�Z��G�$�C�jg|��9I.��&�'�C~�'w�p��ҝ�+�l��Y��@<�js�3��<h_͚����qI49������]�������'��7 t/03�\��J�_w�i��
�x�EVš��,D��$�
��}�!;�-�L\s)��]�
簀��J��э����vLzF����v)%}*C�`��Е�\Ô��:����,q��}9��+�B��Y}�E/��g�!���3� }*���c�xb�y�e��|��٪T �/oֶ���w��wC�R�ry�v�0�x~O^	�u�p�X]�Y���ޑ�G��>��&<*����pƃ�_���ۂ@�;���
QRKIMfy��+O7�9�k�n��}�w�Z�Jۄb�FR�t����X5H��v%����<<�?�.�����xT��ox���j�H���i3l�ҪEK�yi~=��%���UD/X>�����M�ʤe���1CD7�Q��?[�w$�%Y<K������y'#�{��c��o$��F�T�!����t�"�L��Ԫ@��9�L� ��E�tB�o��Z�e��0�fPd,��(Ӝ�'�PZ���A�C*�ԙ3��ɺ��L��<�4�$�z?��%M�������NX�i��S���  �k��o%j���w���J���#U*ʦ�^rA�d���8�����Q]��a�����az�N��ZI�j�%�6w���1�[�X ����ӮϜF���<��F�r��AG�����!
B~��b������P�6G�
H���v�pv����ѣU	x�WƸ6QH
ff/��B����צ�UBwT����]��w+g�.x��E)��x�#��P�����k'2�#-�5�8,6�%32��0�'\*P0"C�����6Bq�D7㥈�M��L�@�WBCt0C�:���@O�%�W5soo䅮�7��A��h�$���$Se5��� a&FhAǠqP����c��S�"9�����R��ڗ=���z�mZ8��I�sf�6�~f�|�1���wM"�r�D�m��� L)9��hݒj���4�*��
.�Ll��Ι��0y���n�`���q��Oh���9L�C��p<p�`3�;m����,�PF���+�]GO���kK�1�-���]Dm�~I�' ]CU�tT����T�@���tɠ;E��{�I��>��6�d�03ꊏg�=�`�(�6��$TO��0�lva�/>�˄Rr?K�b���P�4�w���!��8eq����+����>C��BkQ2a�8 �S���_a��W��=����%Qe���"*��Bw:����ghR�w_���%��(�I1^���R�hs���#�`6;�$�H)�Xܨ��%d����i�D[ \�s�id�S�>=��-|�|�G�g������2� �jE���r�zZEi;����p�
"���
Q�
�}g�g��'Q��8R�e��=�P�IۂF��:h�8�19:�⛃Y76�#[�/�Gv��#7�U��,��{�?����� ���;���"�,��@c�O��#����m1��������}iLI����h[�f�P�aZ�5�6U7��yZ(L���T��������z�9"Q����tld�^�e�@i�խr,/�g�/��D6�i5NfJ<D:/Q+�^�|<�s�d��� 5+1|��p�A�'��%�q	-ƩDԸ�=tY=��]+�q����f�8�6]�N�����ܲ`1]�|ｿ}��L�h[l�!�,�o�\�ܱ�?l����)�ѦS�
m��d�>�n�ah��F����[2�u����uZ#YF.��4'�mXP*A:�iz�y�?�QP� ˩y�j�tdYLV`�zQR���#�%q�=#C���)vXC��ͬ[:�M������޻#�Jnʈ+O�6�A��W��x���1ӛ� ��{��cvJ#�J
�j�p�ڐ�V�dԘ�:)B6���������zk��Rԥ�~s�	k�L����C�e~B�ɛ�y��q:~�;�ѹ3� ����z
g��k��`sסR�Dlk\Ci����iXJۯ���IJ�ZK�S#�ě�7�	ߠ�:����R�����:�@ОTj�~m߆��:^`�����!6���W���yB��S��6�1�*��$�#�?�fCpOZc�(��Y5�x�mW�Ct3Q�aㅥ.͌/V�a��N�ɠ����|^���`#�����h����R�̕�6�k	*���o{��G=��)��}�,ˍ��B{���>c�{h]��?i6EU�@������Q'��m�V����i�cص���Pt�*��O"K����]���F)5'Y� �Ӌ[�=e��o������S��Hͩdk�_]1�(3�*�P��f|,���qK�^�
�Aa]2�^L$��lX�p�"I���gĸ��b����_�TU���do�彅�x^�9N�*ע�T���$����X7��d�YA���V�&�1��MWȕ3���k���k�oɞ�0�"	{�x&�pm���^�%�ZYҚ)]�m	O��,v�ק���#��C��>�֧�̢'5t�7��(��rN,¼��+�q*V�{Z��h^oJ�F�ˉ7lI�(�B����W��Zz'V&�F�
 ��c�g�X@��j8��M$%�q��l�8�D0��) ���d���X�F�	�M�utO���̨���:ѭ���Ф�� �1I�,�2�>5'FB�y�k7�p*��ok[%����Wı��W~�{�u���-_�y���~_�1m��桞jd,��.G���GH���M���x.�dX��P*���[��n�r4�h���`�>�AwZ���3�o�0�n �ƮT*4�I�l�S����XRp�lh��3;[Ss������ʁ�����I5���X�w��οd���4��g*'��Ha��M�0"x��1^������ ���7�޶���'%�������TKݵ��R�Q��h�ސy�c��TQ ��;~��<�՞��2�}�l��iF8�斵�vFS]�+{�]�O3������J�v�t�m�΂Յ�@C4?��L���p�ҭ*[�"�����u��S6S3!��б5�5L�QM���Г��}g'6���������7f��!�$�F=��$.��&`��Z|��S�%A~��z��T&�������4�o��PU�ر�bϡ�ְf�*�LO���[=t�8���G�h\���{�f�M�J�<\1���=�s�W#�&��;纔�w�Y$j�D�PK��G�����5�������xC�2�ڕT�Z��k��=�~w���v~+fM�.�`qMpm�@�ؼ��L�K��N������
�k(��D~��Hm�%��,�n����î���7ۀ���n,��+��D����ӊs�m�
<��%���O��@ ��L�^�e� з��B(2�$�?������y활�Qw��rj.�����m��̫�Џ��_8cў�~0CMRٶI<� :A���f�/t�����+���xk��j��h����J�f|5�I�Ѥ�(QE"i�3���`n>_GEh�;�p��d[C�z�Z�ϥY=5��q[M�sظ�W~����*��AD'�0�R֗.hF2x��Z!��!�tj�]wF P�[��A����&��i`�@�ۼ�����.���v�<�&G�����
/V�Y~�|[>BJ��`�&Fo����Y�%����@
>褶Ϙ�$�`��m&��*����Ң�����3���f�
���#q����y$��F���X2UH�u�L��Dl��1��`<���u� ��F ��L~C��X�5�	��tt�u���3S��Q^���r�Yr�]`���v�	��Lx��+����z(�hW7HV�ow(����)$� yr�$US*� %j������+�SW��Cv��c��3R�;��%��]f�f?0X��t��R�;��C<J�6qb���I�x�%ߕ�q/���Y��h���ג��H�pR?�U6�nl20����Sd��2[}81���q\�s��NN�9���[�$H.{ �*�P2�d��=y��}҄>�a��5�~�=g
(/��G�"�������z�`���C����j�sZk�6�G�Fͥ�;�����Ÿ?L��p�,K����}~_Es�Ҽ�5�ko��L\*?߄9I���>y`g͇�6{�����dհP�Ȟ�&���*���>x�xԐv@X�_�v(�i��-H�	*�0���C���`6��/P�������a��&n�q��2�z4Bq�\vBAFM�߶�^ρ/��9V)SF��F�ѩ�S<�`��/����)���
K��G� ����o˃�ʋ/)Kd�*XI�X�ƴ��c3K�H$�5��
53�nz�>N�𑷱��E���:�nA@B�78��0�'ԗ'��y��Ӳ�v�}�2-�u�K�
D���R�T�#$J�ǃKGr��q�z�V��}�w�q�'�Q����t�r_bB�x�%�T`x� �g��3
kƅ^�c�����AO���{�&���y�X�*"�ס�N�|��E��5���[IIQXD6��E����C�>����,����ʇqų�#sY~o�a�KK��m��@?\�^�WZ� D���z=�v'`��r"//q�V�9��B�4!ߤ.��� M��&����6�1�@��:qV�3{��Ӕ�cA�;��khs�S6.�.����J��,C��.G�%o�QQK��O�l[1����r��{x�m�Ua��L�7�h�����K�]V)����|{n����o|�>���Z	&�G�L�Z�x��\������\ �9�\v�����w��!`=�'�Α�iž9������ǆ��()�&E܄(�N�hr�a:JE�CO�`�gi�`������Dҹ֬���yR@�64���6��ہ�����͓Y� :������5^+[�<Q��N+#�B�`G83��O�`���j���
��ϧ)`�B�&
g��x�#�x.��u�>����?4D�M3O�k�����k��F�e�<�)"PS��S� ,��L8r��~#��_��宾�@�L.|I5��\�aS�̢ϩnj{�,��w��>_CE�t��,/�r�ZŐ���ڵ��JN�#�ܹ]�喏8����_O�r�*��)���������̶��3}�/7%,��������r�|���?��0��{�j��U����R^�׷��z���<:�D�Д�ٛ��4�mݴ �IuF��14ZS�B���=�WU� �ݘ���H��):{��}�B��D����i�q�t� �).F7CA��ɧğ�>�V����+����俅��IV$� �]�4����cT���b+(���Va�_��_&��e�X��O��C�0AIf��r~ļ1�JϙR#J͸���� lת��댹�P_���<6Q�^�����!,��a��"I�L�z,����x:�f�Z������]R>�K���W��-��?��ig6�;"�]RZDk�
��&}�X�L�P_��'�������ʵ��B�����5�1q,6<X�O�:��������)���Qw7\��֜�=6q��l]��"	) �!C�-H��BmV�U�q�#^"$��ze�T��|5č,��"2�;���an�_��O&@�c�݃����=J��;����#��u�=%�3H��r��HNX��M��^���wH�!���:~�n�/�q5���EcX�59�����O�h�/)%�?�d7��~�Z�w|V1|���zP�M7�X�4r���T����%A�.r '��h�X��f�򈱀����*��Rw4���N�}ז����^3E��aW��;X�{�a9��-j.o!��������lx%�V	c�V��ټ�-�34C��`�^תXʿ��h�LO*�O��.��0M�$�ȉ�Le�#3�2Ǝz��aj��ljֈ��N���"���LCH�x�)�;�$oD�!9DZY�4ܵ��������)]P��!�Z��]���(b=iy�8�l���Lk݅;0�����Δܒ���:0�8 �3�P��\!ɫ� Ŀ?�P�db���G���|���>@F@V)�����$����QEh��I3ܛ�ƃv$D�贑�S*3�ͨ�x�+����4q^q]�f0��)��>�r痷�����BC<�����o���=:v�޺��LԷ0ރ���Zk��SY���� ���=�F�k���܂2�e=*	��^upng�p��׾�58'�E��Ny���E�i��\�g\�Y�.*H6���EB�Q	�S���9�V���_�� b�m���Xo��:@��Zv��/f]OjcCe|�j�'�x���ő� p$��(lM�{�r�I��UY�1�W]܃#���}��N*8�{�� ���@�z4"���1����n>LN8���-IQ�z\[4}*�@Iqk�a���H���9�Oq�c�(�����,c L.�g N��N(�H�ԉ��-�������6��Х`� ��$��.rj2�)�����?Wa^F��T�~b��>7����v)$�����,%J���{l����
��H\��SGF��<��<��=����p���o�]�~K���/�L������y(��WC�\���+���IP�k����З�J�C#�j
�a���Q�`/��H��Ka�t�I�Y.��n,��|��8]�_�­��U���SV�26��T�]��DK�C��M��nڶ4K�8h�"e}5؉Ѝ��#�B8zc��L���]M�� Ֆ-( �-Y��8jN?�݀E��,Vjj���0���q�*�.*�E���&�)��k�e�|���%��_��m뽼G�{�_D�F|(�yU�����l��} �4��������$��T#\�W��P=f0k��PG��~~\5,h��y����9y�w�D�p��BkdnE9� ��`��R����v5�l��F5�.����,���K��o�_%���]N��Ds�	S`O#hͩ�,��Xf*�sY��0-�saߙ��Z�}�hT���_���2,�u��[|7���I�[`혘������ 'Ď�����C]&p�Hʌ��T��t�0�'��!QGġ�8�7ٖA1��'M�K�A�ޫ,�����=�{���G�ƪ۶��	�=���S�d���편
�*�xW�2sY�.�� �*�5a=�/EZ3h��'�����?�]��!�A�ƕ��շJ|�:B�UpX�Ev�h�'P4
ښ�+�l�85�d<����b���y��iJ� 2D.�Y�r`�S��Z �Z��(�I�1��%�k 2��
�'��z�v������>Rdp�-R	���R�,XX����r�.z�2\t���D@}IW#�QV@u�奕,%Ht�� ��,![\a����}�/�&�.��3�0�.>{��bQ� QBt�%p��-B�q�ЏﮋB%�!��M�N{N����ssTG�;�{(�����7 �_@ֿ����n�?10�"��6;��/p���q�� ��Ifo黲� �����j���{.1�Va�x����W�H�P
0��c�o�/q�w�R2@�:á��T,o%���-��D��g����Y$�V�MY	�*�a;�C���]ƺ��賣���hs��ή�6	�u�bt3Vm���a/ ��?�NꔕE�O"?�A�Txnlb�?�a*���2�~K�@Ry�CՕ�����sD3cܕH/aw�]�\ c�_��P��ej*D�s]��Rb��ݩ��`��gܑ]9`Sψȷ��C� ��=�P�)�c���\�,.����sa}��U�>�Z��B	��$�cp�h�_'�n-�]U�%�����t��G�uc=�a#�-�	�qD0�E�p>���}C1�sN+_p�����_ԙ��&��W��F�V:���"����U<j��؟��/�I��	fU����v�t����Ό���X�P��ڱ��V-��ư��݄۪�:����jF� ���o�"�'"pZ��V�[$f?���U�UX���#��`{��S��AL�ԫ�|*)�>>�&e<� �b.�@�VJ�	�|�A��I�2����� ɺ*�n���eJ��ԝ~ Gmg���.�g�㒆nh��n��>o,�6?�� �.\5���|� FY�3M߇�\P�J�e��&Z��h���?�2m]��ː����V�f<#7tX�|lDEW3�lܒ�/����C;�
�J��̑ԕ7���g@)�6�#f��D�bk���d��^��AWۭ��ݼa���mw$���V �$"O��^'� {P��;/�x��F�R�W�m�_q�YnP�8���V��p��L�Ma!N�#&�4ѐ��S�j��cw� �aܜ�_�VI�q�rw9Y�H'b�����n�Kx."����;���B{�x"�[O�����N�0-؊��+�A��[�1��1{�9���o�!I��"칡��3Sم���J��GT�
s&�b�pS������}B;��m� `S�!myО,�Է��Ӣ������f�k�3��c9�@��c�Hݡ)-R���-�my��m�{ˋu��	,��D�%,�iw��2E��z5r����e+z�.C���%ȸ��k��Q�h��H	ɖ>�f%Sr��x�B�+kZ�H��N� 4��f�\���&���hf6���Ly�3�|p��𶐇ΓY�g)��m)ݧ�H�%�x�1���x��*Ml�w�43��՚	�^�4������戕�V�J��C��s�k�&��Q��n���#�Yu�i������u[�[K�%4���a� 	�$��T��g��9�iE�`���q��xR��m�:ڻ�f�#���0�q�< ���d����"�knH�bj�O�}4��q����]��L�z�-B��/$3 �� }&���1l��dFX�Q,��+b���|#T;@`�`x͛��Y�e��C��<�V����ʇ�nu������P!�g��|������������o e G�#戞��Mw"��l�B~�v�n	�t'��B��i��� j%?�����M�9u4T;)���ۘ6X	�j�ۓ+����'-�p��ٞ��l&XH��M0���hN獣8!B������BwUy�A�3D�3�ɄP^�v��N��f`�t�,�+���om�׉O�
�~�ςU�=����^=�����ϻ�|�y��;r�3bo/��Qu�����=k,���&��룡]7h�C�'neՑ'�}=!��ՄZ��5!��?0�Jtx�pAb@0a>_��I{����/
��p4iXn�� �ȣ�CJ8��
�U=����RM0l�ZۣT���W믐�I�d(�%h%w�+�<s��+̕)���+-o�6��ZɹE��U6�{���i5F�P)���W�T�Z;|�'�),��z�ۿz�N��b�[梗r#��,�̪C�E��w��ۥXB�h��T�"��f����{yuᘢ������'b���{���	�{��%��rz��-C�q�c�J�
��ۣ�w�h�k�TO�_mı����B�~9L�4jLޅ$���t�<�]6W$��%��#PBӋ�I�R��Q��[J�����.�U�KNm�c���=��G;�&5����A��NS8�kF���<�w�"��;�t�+O�[���O|��#eZF)=�PE���oV���l(��� �I�S�s���X�h[�c��5��#�tc�p/���M����4,n�P�Ѵ�N%Y�.,��za'�� �q o��pr�S0m�7�6���uXnp�%=��-�T�d�_���V���c�I���2Q����(�?eV�S0�nd��UC�[��?g2��5Iɋ/S$�y�e&���}�6i���JO����q*�
�a�&#�D�˯1)��xi���­���xP��)�e7�H��Ma��9�Fw��ȨXt,��>�r�$�����ia/�v���?��X���@�Zl�a��5cjC�ú:��I[/ᴆ����%Y�FPVb�
Qa�ﰋ}���ߗ֡��]���PT��������B�3�ʎ��K}�,$�$���j��յ%�?���)�ސ�Q���<.�*��:��][D����B��Bd�`jX0��AF�g�]˗Fy;.˽ѱ��G��ŷ'o��5�EȬk���E���t�w^�.�L~A��:����?�N�'�w�n�ZN��/@�d#^�l�+*aG�E�����rK1��[.�͏��aZ�r����Q#c�/�Km�|@��'�L��Tb ��� ,}^���>�F\;9ԡ��,2�o��Q<�R�2{d�JH�N��`ŇL�X��aH�M;��D�T�wu���[���OJ X���6����/����[b�1{�s`TUvs��D��S��:�T�p�d��3č�C^b����8��[�ɢ���,��(Ř�r7hͤ���Wr�Q��;h+�U�g2��?���
{8r<>�r���ݫ�*�r$$�a`���q����~Ǩ0����k��8�3S=97��;|-�e��k}@��q�t$��v�@�T�|9+�IC��y��ieWu�#d8�W���J�q<2nYB��0f[��(X�Ũ�C����,K��Jc� �<#-��,k����G��v�+lG'QL�C�"R�uB+�rN�t�n�R�㐞Mv�[��e�V�`������M�p��"���k��Op�� �����"�V��8>2h,�/�泠���I�������6�L�K�n���{�E�=}(�TX��L�5������9u�vK�X
W�σh����ż|���|�<З�v����D�c�;P��6��*S�lc7�$"���]0��E�_B9����;j__���[��a�]_v�ђ�Gf�$�Ƙq��#�� �.��xS�#�b�ԵE�d��4��4-�֘���jw�W���3�3��ch�j�"�*�{_����`�:�{�{��h6��Ϳc�t��[�`N���C2�����+x���z�_²�4J'V��${1!��&�B2�[n<�М��͏N�̍;Fb�7�E��k����QE��y��I���6_f�`�+f�"����}�c��H��|n���>��'K8�,��]�-��y����
��ZGI^�q��+�;Z�ÒVa���u�D�&Q����ʣfF%�������Мt5BU$��`?G�Eܚ��𴞶/>`r�F cG#�����R^�38\v��#)�(���m�.1���~R� �t�Ph�!�h%-�K�t�� v�A�N��m������v}	?kej#�[4�.0*pq�a8G�B�u-<�#��E��#(3��Cv�D�s�P�(�E�<���PIs������g�tTt�Ʊ�5��`�g�	H����Q�B�m�D���g�*�_c�"E����p[$��y��	��L��|/B�#AnUg��>$��|H'�żu_�O��W�K��MG����Ð�g$�%R���fI��o�V�5��v�	��)�P����;
T�42{���0��oJn��3���T��TH�d k��0�؏��>����`6t3`�3�yo�~�fEtBEI���	Ɇ� z�SPk̑q��Ac��{�-S�b
� �w�_��?S�'�f��5ϱ"�ǋT�_}y�8�����I"��ih;H��5��M��Ȋ&��'�嚃X��<�17~�Ne���;��	qD3��r�$h<(���ZUyI���o��I:������Jr� ����e�yߊr���$��;� u0=�NE�g�R��J r<��_$Gg��#��B7����"��2�Ph�l�0�>�֞�4�
���_��%;��1�Ò>����fg�С�<�
��νZ��R�}��VtZ�K-{x�)��;
J��x�IwT3��5`"�����(d�p*�h-��3Sa'�P���=M�W�8R�`u���+˹r�Ѷ>%���	�_�����<T��랈'�d�B��61<��Hj?
�Thq`Lq�V��ǫ\m���BZPZO_u��� n>�C��x��j�5��2�l�������D��< >F��W����b�:�����]��' ��Ѭ+ȔB^�Tv	��F3�Sz�/��e�C�>g��K�F|z�/�%9�ҋ����{��ߑ�Cv�9�t�~����5'i"�0���(~�T����3�OxG�5DzĹ�ݯ�%�/���A�B�5Ƴiby#s�[�%���M֡`Y��a�^q�@���_�g�$����f���/�,IH9�s1=�աZE�M��rw�QY�k ����p�Z�9}�:nOP�uH 9�
���]��vE?Cal��	�Bp���٭d���N�LBc�pQd��Ӷd���-��*彅G�)��C/��)b8OU�0���sCՒ��E���hsDI�mL�ϐK:�@�\���8�7�N����`&�gR�ϱsm~�5�+������e�v׋m���c���c�UL�������ﺺ.��)(e����J��ʸ=o��$��恊�&�Yr2�Ըi�ʜx�"I��%n\�
ɕ���6B����l��S��'͉)f;�w�(�����w�UH����^@M�uE��a�� 5&�CB�k�b"S�����k�A�Fی��wn�
��Z ld�JM�3�Y(͛��KOf��c|�t�NM'(��w�W�����X����� ;�%���{/7�<s�ҽ� �Ex@��4{��l���w��{��.���}I�'���`}����OkEi������������$m�bױ�f���Qyx+c}�O����X�>X��O❃��bRi�A�)�M����������H���I���w+f+�����O��=�=���<�`���a�b��S���Pr�\�;S�<��!%�6Q4��鍰��t��xA���.&	 ��t�PLv��±��l�Y�g�~�7}es�dk.��`�:]3[H	&���L�����Ϛs_����(��^%�p����K��Yסom�+��Bqg|�ߔ�SU�a�0���w��#(��UiK�8�ލ�v@jQ�Z{GS�e��׀K����g_c>��;�bVb���5�3���V*���b|����#%��WC��$:I�?���j�3�4ԏZ�<]�X%t����R	�0!��;j�������=�ѽ[[R�ae��W�E��=�yd76Σ�H�c��^�A$z�r���.�܊�5���[�I4w�nu�?�	vM�,��PЁ�Ʊ�?Ag��@<v9^1��D$뛜=���$�8[>8�y���Gd���XIwc�.���η@�2���M���^_�M�͆V
��n�:]Bq�7������B�ww������)U��hD��d��Q�O�@E�/�u���i1:Ht,#���f�m��1%B���xmBa�{����X+8��l֬���Wb�����٩K[A �L�&�8�
�=>���\{���(��,��(,���$��mG��x�'kZ�)e�R�F�4�e���E����u�4���=�
���$�E=PC�Z`|����M�ʌn�bLy������g���$L���"X��D�Ri�9�Mge�j�����'N6i=M�z�L�� �	+Z))�OBn��x �J��1_��]�4������]S/���V��$����m�� �5��?ϯ���VW���Y%�J��_B2?i-�I��]��o��L�xm��P����;��l��y�:}Ff�IZ aDJ�|OnN ;�����T��Ap���E����Ww=�"I��E������|�cr�{�z(V�I�هv=�B�%a�SK�i�Vv)yO��@����p�>.��Ll��r��律R��oye(`U��#�=�%%�N�$cGS�( F�X�����"t�1�*� �=c��(���zɀl�Ҋ��jE Ū�w��4�}����#+͞՜�	%�aáL���r���P��-(Y�!�U[]���8W@�K�E!���V�'�����8���ж����ХT�i� �-�N�G_�Dg"��)b_�'ap'� t<�O����I�u�D7�V�Sά��Y>�7�Q���6���>�<���0�,�5���1}	�<���t>�J�\'�W�>�j5�%��}�|y����%&^$S��.��˱���"&p�t�N��v��M�ec��,�c������0j`epY���i�ʡ�xD������������* 
��!�����hh���-�vs@Е��h���;� v�w%6���9�1��
�@Z@Y��{+�9k�A�����u�^�&�UQX�z��`\���3�ԍ��!��\���i���2;%�)1'�wX�
պ�1O����2Z�����!g9��w�V�iu9��[�R�;��F�����Y�h�iq ���-�$\�j����"�b��"����!�g����:��q�*��|���d[㷕���T��}к�?GS݌3��/�n"E {��(�+� ��i(�\շ��'&ڬ�M���Q	�3:�ź�����!k�ٺ��J�ZJˍ?{�Ȋ��s$_�Q��YႚH֊��|���[�]�݊�W�`�-^K����ϔ�J��
�՛% ߬E�+��Խ�Z~]��ͨ���}ս�aX��Us@E"Y=xHw�nQ>��w2\���G�T) ����?�A�)<�VV<=��+j�#���	����\У�{�"lյ��P�oG�8x�GH�$R9A�ȝ�8VF�j\J�tށD�c���m�^��i��q����;:�]�/��Y�V�*Xx�cD�2��W@�%��Dj{�Zj�_� �ة-r:o�8����W�L�ǘ�&�9�p�b�<)]�ض�主��5qL��SL�.��?s%��
�иj������N��s�{ϖ	��+�?F�\���3$���{?��ǻ�*�sI�i�h@�#g([��dyc ��֟H�y�Q��|K��d2d	3��%=.�S?UK>�����ПL #��6�W����TS��G@�u�R�X9�W	�zƖ`C5|�pPk��L���jD��d�4П��AA��Q�.���,a��O��H:��VI<�h
�47�#Yw����M�-C����R�l|�S����Z��И׼k��li�7��)5�zQ��F���5�LM�UWg<�
�t��D�<kd���	�:lKIY�Y�~KD	cYo�%4��Ow���j���=}��U�1M>��ρ�[�=�	v�B�6�v�;����E�u�v�ͮ�T��ѣ�u�k�Y<:�� �7^yC�q_���[S���:^�:��-�df�|7���~���\W�˳�#[�Kl�%��Z��tj>�Ԣ�mܻ���b��J᫜g���G��?�[�V�����f��%��R����2�.��)��՞�p}��i�o�����{B��=�8����%��Lk�y�Jv"7����WK�Чc�-Ĥ' �вYiQk�h'�CR�b�m���۠�1��>�.�>��������(�M�	�qHp�=Q+�2)�{�j1!��`z��fT�ƶ��2/ch�ΩV�tgtIV<��D��{����c��@��o��QtYx���B�>&Zm�.Ǹ����f�$bRm��mw�B��h'ͤ�W�Z�+�V.W�L�g�ޱjS90��@gʅ�!WǠ$�ϼ�`��,�0>f�ܻض=6�!ӅTDI$�3���# {tm' �˫B�&�
-��:��A�y˲���h#`��JU3(<��@�#�
�m�V�Ɖ&����?yb8�M}�b2M)�w�z�<���:��dW2�r�����(#���5b��Lcr�ce�w��\u]6�N�)�����N(4���݃�Q�'G����?E��\�!�└z���Oi���	v��Tf������ Z��״B�G�~�ׁ��\�r��#�Gmv�>G��<Z"�0#"�&L�O�����n�%�"+ٖ�@5)/�z�.�tG���=:����8wt��SX�\�m�����8�|�S��I�f�0iS�@/��>���)&3�E�;��4��)�;������	���}k��'�n܅��d"
X�@oV��)����e��]ly^�~� ���,p���'��څP-��ۉ@�ѫs�`����]E=���S�KQH7�-ŉŶ-�R��w�_��*�j_ ���a���A`+��ɲ_�������ny�;(Ű��k�''��_yI�
o4�貒ݗ��d��h΂Ű�en\Bo�{�WZ�+�\Tԛ����P�̽7e)�~8�D��rvQ��i7��ŋ��HN��4���peָD��?
��}��V������*H�"J\s����$-������"��N��X�"Yv?�_��y���n"�]e��ҝ�>r�fm���4����r[5G`�ʽ��h'u���ug��*+Ն�x����.v�1�I��s��E;��O�j_�b�`���{h=)
�M��|M�[n
Dؘ�c�cOK����l��5��W3v�DO�y�Uxܒ�Gi�(5��'�pHk6Dߗo��;������^r�3�|����z�;F�����ڄ'.^�
I>��N�$�G����_�=G��Z1c�sB��j+�/v4�*�6�1c��aG�k�T��:�^Xg��]OJ/��B�l��5_�HU��bzY��K!d���;�+�[�J2[Z<�P}��˴K�F�.����L����������uͥ����d;�Ri|˓ޕg�bZ���gQ�3!�}H�Z>��=�����5����l7��T���u0��]o^��8פ����p�ˢ0nWRT��FR
r�.>8��-w�A"
�/�}{K��Q�)�uW}��%<�]ϰ��K&.Ѧ��V#���68�<TW�?�#IA���%��(�2����sy�R8�����ԙ�"����m+��vf���?�<͛�wD$g��������*�}?�g�����P��)�g���B>�5k4mk��I��fUr�6��Y�T�=[ZԖ�1��6 �������b ���knQ��+��et��\�����(E~��.�/k����0^T��jI/
{]���hhl4U�X�O!��X��A9�弨c?U���ܼ[9�YQQ�����P��E����n0�ŨL���$���4s"��@iw��`�P��ڝ��}�\���#��y���+���Z���?;w��� ��'�:χH܇59���������y���55�E�!9��`�4����/���2sEy�k����?�n�8U�*���u/�{��ܨ&zmj ��g�(bk�q�\䍺>�4���D�f(&�4�d�-Ag�}��0��e��J_7$�/y����ռOX�7��\"[V>_D{X�2+����ꛐ<�%3%]��vlrx�·8�u�A�Ќ�	&�n��*�l�$��� ��}Jr�]Hdm��?�˝��8ᡚb˶�^�pD�*��rC�~WED� m'd���Y)�yN��� �ec�O4|u�y&�7�x�,m8	HE��b]�
�|'��p��l�y�T���nlO������p�uoa��Sm�{�m	;��l�1��h5�Iwk�	qp���U_fz�a-�(�6�OW���!\ې��%�P���+�!��P�Gzٳ��ვ�Lǯ	�hk�i��U�l���O�}��
���7B��ຼ�/�^OA���O���
O����>��eL��݆s����tPG�^�	V�V�AH��a���?��?�7�zq��� ����Ʀ��7�M�Y�N�7��e�_�U��u����>�Z�S�C
�Bsj�.-��i�	r먡Җ��Y�c�e��δ2C�a�qj/��*�< v�����<�&\k����������� ���e'2��O��%���R�=w��M|�,W�t!�aZU����Fc�peo�sOQ"b3��Z'������N8�شZ}z��P^���2?�M	M=_Z�}�}�H�ɏ]&(27z3+=1�(gB�70��@����T��jv�j\���ĩ���F��aG����{^h�' �ު��7��E^ڄ�q����clC�;�RP��n���]x��<A��I���R�bq�Y^v�о�Ǭ$��Օ�\_���|խV��&!�랖CqI�%�Yf`�E/%���5�+�M���T{)��Р�u�d>��64Rф�k�X8(�OLA�o*�ɞ��|5~_�Hb=���3����Gs���l��厘�F�Ϡ�dC��,�!�������;����X�kUU���`���Ӧ1��L����#��R��x�
šWE�)	�4��%E/IP�l^0bz�3^Bh|w������� aD�@L�f��߹��y���R����Y@�j��|��u����)��>Ǫ��9$~ܔǀ"�R��ڇ-�kbǾ:�"��i�m6m?�#8�]��7��9��O}����R@���P��6����Q�2�b�̋���-cT�|�1���V-L�	�g��+<�h[oc���|�����h�k*���S҉>%G`g�D��eO�!9�GǇ����mgz���s_���)ޒϼ�~j,Qv��O��R>��?�s��Jp��n`m6�S4JT��o���'��NǦ���`#�a��W��2V�9�sc���w���O-�� ��+�ς��7�����#���м�a�a-�K����.Q��OB�*�s�t ��l'd��7BK�A���r��@t�.)w��i`��z�����3��4g��+�����v�V���;�'���*#����3ˠS�]j�Wb�ˍ&�N+af�U>j6����)��!78��tiXv�o���qNٞ�k��C6&d &��SC]�z�22]	o������J�z���t��k�:��Iv��,w���1�>�#!�^fւ��mh>O�s�-�ǭWPI���2�/�2��-R'm�Ğ�PWة v(����2�a�і����۱k�2��n�j5���]��s�.�DAgL2~K�k�49ae�_Ы����
aF�����)@���r�	0^�x��E�<���[_	?��,�,v�j�o��3@H3_�k�蠑!����zA��׮aב$�Ο�Y�R������o���ir�C�L�ı�q��:I.���ٚv�������~�99�#y��9�o��S|Ys#�N_�432�6eg?�����/uXb�5�Q_3�{x��כ�)�f�����>UQ�JSp��G�g���'�3��[+'[�])k�tl6���,�� �j)3/�F�������ԑ$"��:ZJ)�v=���{;��
z�C�H-�t5 �=�E��V��X�y9��\y-T��/�@��Jy��[���:�>���C�S�$��%�8*��������U����B�θ�6��eO9'���D�/���5�%������˃���R�D��{�7j�]�����۠(�M����Q�I&X/��,�'�:P/��`D9���?3����ڶ$��ZC��*�w�ϺN��Z�y?��=1����2��ޭ���xbR������=~B��~\���Uz	��A� ��m���X�cj�D�/��|�v�R&�=0_a/�QR��~#%6�p�C��,�� �h�A���u�h'@=2�$�T�����܆�g�	O��=��f@UC&ed�c��-𽗄U���ĭoU�\�!������ru��:敕�MLM�`�/�%��i�_�¸���9%���y������4���S�;)=A���3���bc�@��'+�d�9��^�O�3v=dB4͘��=�(�Z���6ˤ�vWe� ���:�� M��1��Իnu*(F���q7J��ڊQ��g��@��h5La����_�G�Gh�>
(�[V�%R�@�<��}���3�A[R<>S��v&������&7i�7�rt�ghEZ^{�!��/�"�>���M�B�B�1�� �!�gPyu����w���D�M���@1���6����.���B���)~a�
&J��1?����z�-ri��^ZGlx?��M��?#H8�m��o;X����ʠջ�������XU��k3��N%f�i{�����]?��j�����c�\<��l��4t��>�M����c�W���m��Ǐ������=2��}N$$AU���j����!m�Y��|Z��	��t���Xo����W{o��?:TsD�o_P��9lH����'�������SL�ysAbќ�����<�}��I6��u���5�^2�mh�g�9����>���/��i��b�����#�44t�=�$�V�CA7��L�:�^e<{�4�~���c�/?���+�/�Փ�e�[����HjU*K����DgoBIRNK�mi=P�Z�#��
�s�{I�_ћr%�-��Ϫ�C5�5��l�!�z�=�����r��s,�7W��ze�����>&^9�C��꫙��_=��[(m T:�y���9�8����-C�Im��0&���(�3aWp���)��z'x�1Fs,�N���oGB\��v$���������k��Z�����pJ�����2�}��Ч1f����ꐩ�H����^�vr�`轚)�G�{��=d⵫���,�:)���� �	PwS�	�n�;�����ꗔ 5x�ǴWm�Uߔ��kX/C��it��_�^�P՝Yޣ�"�7]H7�Zࠫ��3T��H���޹/X$Z��W�j|N�歭�t����7��D��2k���q�m8���r���D�q�@*\D�S��3�$"mĊc��AO댠@(|�vNo��X2<�Zd�6�������ohbF�Hz�� ��m��Y�z���L;=�s�k�r�b�O�����ub�]�w�~2���9S3A�[N#�{.�L�(,�8���2��e/�/��+�w��<v|*�����!	�H5*H�:1�Cbnba5���#�Z��z�/����^rh��B;�)T�Y�5㝇*	S;N�AF4���`��ɻ��*�׿�!�N����6o��N��V��N%�����[R��,�ɖ�f:2���O�]����S�ڣ� �M�p�sGV=����������pXZ�Zݫy �'gv�aR1\kھ���E�t��:�X`'�%2*�B�?���DX����߄���u~����$a�Q|��R��3S�5�p؛>����4"NA�qgL�Im�G�����d"J���%v"mY�яU�!u�ѸJH_��Ƽjfa�@�vX�:N���j�S����륨���)P�h���|�ju�%���@j@�v����A�j��j �2׼+&G#�ecXr[�Z2�NϜ�o��P�AZ�hi�l�0�+��FtJ[����\S*Ij��w��Z���;�ky��UxS}���$R���3��R� '���A�'-�=9@SK�i��P�4�qX��{�����-8�)�J���Xԩ���}�²I%)1L�� U(>�<��=\sD��r�A���8N���]�*�!����]����H��hI�Lw��؀"��p@c�&�.�J�+��{��j�P���:��y��J�'�yT7�}gO��=M�5���PfJ9�����H�E .�ob.���Y� YL��A�T4�8z +aZ��(�4Ǧ�X|�%)����d�=����T��^�dV/�dZ�q.���@ߕ�C)F�A~kl��R�����.y$ȳ�O�	��;j���\2��2�ɬ%���Q�;���uT�^��oש��;_���Ŕ%`2Hz�|PW�m٩��G�^�-�b9 cx{*tK����d�XE2�8Ѱ_��Gc�Є�����ӎ��vC�Q%�qvTkV�Nש�!gי@V�*p (L���DIUP�|���@#��V������(' H��08952*�@W������Iŧ;`��]K6ς4U
�C��z��,��Ɔ�P,8������`����3��}�ˈh��0������	��Ȩ���N�e`;0��K6�9���궑Q"���.]V���E�R;3qs�V ~Ă���2ƴ���A�,���h\Q�������J����|�ֲ�l �xZl�I��^��m�6���� �r*O
���9�� �?4���/�e�y�ƶ,�6���9,]���]���9����	�^��Ԉ��8-�:^U��8C��奛Od��[HO���r��1��5x���'����'�)�M�{�YD:����o��
��+���<'஢�����j�Q�<��^���گ尩<s����������>�����}�������	�u��� T}��aO�!�[���(bL�_5�B�UD��B��9[Y,0&��.� ��V�Pf1���@������P�Q*FP�Rm�?6�WQc�9#gu*N�7�����d�X�����
�#l�o�ۮi�ʿ�6���$/(9�G�ǥ����+����ɃL"��T��0Yٕ�¦��kI�;Gl䂊�ԈȀ�+̜A�!��<�*��$"�� ��?k�w�d��|�����@�S��}3J#K���_6^,y��f$�����(����s��-���1�u�	�k���K1&�v�,�J)�8�R��N��;�6r�P�����9�#��3~�;��[�R���b^�;�� |�D"%��^|tl�F5C��z��,a��2ķ,��A4�k�����Eg�I�ǁ(�2��n�Ϣ��,�Fѩ7�5R�0DZVB�Ï��@����<�#ӛn<��#X�E��=��n}M�����!��V��+VgE�h�͢B~��6�|���d�R�妉�"]���5S�d������̟��ץj�wq)�PJU�7%��܏�s����G���6�X�A��R��&�>}&�կ%�U��0��i=_.����YOے;�S�F�U�^��c;�f_�iՄ�H�-2KtF���bO7�ܽ=$���f`�A�o��^$}������Y�.�\u�gX�g㛨p]�5�c�k�W�Y��8f�����Ʋ�� 4���[L�9�e�����6ކK��Ϳ�TC�|���C��~��y'c�R��T�L���+bO�7�^�����N'/La�J��k#�
j�LD����Ҫ�_׵�F;�0�������/y���?��m�5j��+��y�i��bW9��+�p�J{����4��j6�R�=�vi��A�6b%�l/G���B�Ҩ���"��Ch��C��������/��>�#W=^�jv��1)2W)�C��� ��.܌��+���p�AL*�5�Q=&V��S��\]ʙ+���$#�>�̰��,35���!PP;��Aw��	��1-A�FJI��kV�fc<1A�j�r�ꓼ�f�|�q��v�cC�4�w�b�}���2�STʢ9�tb�\��)���l�}�Ȑ�䴟��t89��P�	�8K�k`d��&)g���[�V1~㗦�j�CF���j�\VC��q�����0�Y	0���+� �SJ.L7�	�e,��߬�7
���7��iS�����%o4ɿ[��x����:���R��a��T���aڟ�Q� ~���L����cL�:B��\i�խ�\)6��Cd1$Ci�����9٫�M�jy_Tr����r�n��5O8<��J� Ұy�%��e��a9���T/e���t���Y/���2�MA�FO���<`3=���p2�ɵ�y��|�|�m���&==�x�su�Ӹ��=��\��]��,�xG$���J�I�x-�������-fa�\�[.���U�u;)���|��u��7(j�)wo_Hȿo��z��_T�,H{J>�3k�1\$��L� �=N����}ِ��/�Q%X}vX���J4������O�W<�ܴM<��{��n��}a��I�7�Z�{��&.��.e	�k�� �@n���U��'�PJv[1J$5A��5LH]���|?]O����F��Fy���j��&ى�ds�*\�z���2s�����PK��.ы�j��2�F�$э�^d�d#/G<@��VT��&8���3^�E����n�N?�5�6�2=O��2Q:	QVK++���`�;_>�Wp-y�xi�(e��&p���ɓ;���D�/� P�,wx��~U���c��d��Ws-�Յo��EPj��h�7�*�F\ @�\ ɼ�/I]�����!�k�/�侎�C7:�	�+<�9(�L���3F����1�_ ̐��{�mV��/u��cepR�А��"�S����("1k8�NzʦF���Vuy��1^\Q1W=�k,����ϗ�m���X!�zA0���w*)��J�ͧ�����]j-�g���s�yLǓ�c_�.��0Nya6����xB��3�N���wc2 Lmb��}���U&M�_��� �"A0��x,OE�q�HB
�>J٬��r&q^��H�$i�&㙍dt�<���?Y�G���C�8�t��-�����TjlxƬ�����D��#�o!��=����k�BG��I�%��*
���f;���
�I�aa��՜�'�]�=\0�#��5Ql�;Z���W9~�4݂�z��.{�K�Z�Sz{Ta�\ï�B&��n����mxly<�Eև��;�@�&�(~�?5��jూ5~� B����~^k��ɹa�H���L�[����Iu��$p��������͖k���;%�3���$�u� �J�	���x���N�����D��$|9��[IU�o��֋�'��/ῳI���t|,�ʜ,�m"��>D6A^Qw�,mT٫XIDbЌ>�ƪ�q�S����,c���4��ҁ6���;Ҷ��(ZT';8�qa�ق�.j�~��(�@��!V�Ҵrޥ��KIh��w�o+g]4�	8AM���9�ד:XY���/�?�����v��m�Ð �h�)��Q�	/�~����ȋJtj�Y}��	�M���R�uh�7���<�;���fB�3R�C�l@.����Ku+�8���$'ݠ��=4U�� �W3KV��tS���k�D͐� �.�V�FI�v|dA����,�ཙ��wl�d`[{ٛ�g�~��褾4V�"*�x��G�m����c�4���R�I�h* 08(GV��b��j���صH�Ng1�����ʩFA�Sm1��g��|�
漿����u�P�"�/$tBM� ��rҟݔo.�_�u�!T���ٚ�����@D�"#��|�_���K�X3��kS:6FH�c��-[]W��]n{�d�	B����թk���\�k;��'��3)��G�`���C�hlX��
�UB�ę�h1�
!�C��_�}ި�{�WKW��z�ځh�:f ��1�"e
����pSSQ=V�$�KI�g-���s������9oI�m��5�kqCF���]oa���Nװ�bT�MF���Tz�Mn��+�����f��9�?�E��n�јz�^�V\��yV��@������ �i��y�b��	�~U=eO�"���v�A�P��w�uy���4����+r$��A��:�Ca"�$���Yɳ���58^&����ƦU��q2i(&����E�装5���-^�r�[W1�����!���B��j�Gr�6��Q�*��I��"�m�^ɓ��m��c!T%,��%��1�u����v�cܨ�u¡Rw��l�EN��$���d+A3�a��~����R�~�"�^_B��]g�Vk�Uַ:�h��c����y��k$��a?�ƞ}��0k�E-D=i� -!��=�ލ���:�c�)PYrA�N$L.fC��IA����5hv 5*���Q����b�$�4�g�K�	oh����ͯ���I4�9�e�Vb	 ��F�(ѥپB|D��E��1���_�h�z���H�UH�����9#5���C�Z��Q��V�
�����ƌg�ˌ������$���A����bcR1�Uyݜ���S��K��1�^��6t�Gve.�|�j2/��$���|yh��R;ϥUL��p�o��8{�K�����d>����zt9�[Z�f����%��0��KR�ٸ9�\�ů�Ϩ�l\���|�!�isE\��;K�s�.���R^�4?D�Ȳ�[�}c�e,P��5<�f�;c>v������$�d�'O{$������� `��^d���;5��&	,�Ç��oFקI�k����+b�QE�7D�)2X�kKϙ��h�݈�	���w��Zl�㴺��~���̨�0���
p�����;�Z�c��WV�C�Gh۾A��N�E5����6y=Jַ�Hb��G`K��T�D8(������2u)���X���`��u���E��#�`�Q�&@3���w���� �y��Ŧi�8�m~�\ΠU,s,}DvGܙ�t�n{-�(�׎�D��1��"�O�l1H��. ^sǤ�߄�w����+�ش�0���8� 8_ā�X�-�ca�a��/������|�瘚�p��?w?�P�`�n̀W¹d�T8�����˞1	G���'�����|\X�+nu4'n]dizC�qC��֤��~ܙ�?�	�H�?�;'ڱ1�A2$�c��)6���޶~�2N<_t�)l+ԃ�R�ͼ>p���7��_���n�P�c�U(?���3E�t��v���S���Dngx�Kب�dz XY���L%%����h������^������q�Ά����(�k�� ��?�q4�ڠ�Z�v⓹�8Mԥ��g�N�}l��r�P��$/{�RQ=,����lU�\0�]��)�bI�؈�l��4WI�*�x[(��ٳ�#P� �rT���=�+��;~$w����Ɋ>���Ғ���3x8��݉ �7��h����O�ȉYF�r`�A�-r��_O��f�s���ZN���z*��D��A�R'aQ!Sb�3{s�U�țR�J�%�}}ם���SS[3���~TAm��X���[	�;YG�б)Y)�p����WwN�\A��:��$d%p��l�l�����r�ף'|����s���,��c���{�'�c~o�v_@�ĲR#x�T�Ѭ����lrF8�rRj���ͲsM�Gʣ�i����[B$���2Gk:�����MI��ܝ���,3�M���W���+^-���G�XBO����+�n$ �Ν���|�e�)�O����o�8Z�<���r�$0�P	��C���G�u����	���e,d[r!�+$�j�qC���i�C�Ui�ʙT�r�H�/[.���H�_Z����j��]���7x����cI{ь��;�j*p�I�ď�$9da���OM��h|-2�8����h�n�EA,�(Vr��'S�/�[������
Ə�E
zvr��m�io�h�g��S�&oq������fҀOY|Z~HUX~��юEK����{�bd�&W�
����
N�F;�|��qP��/W-=��f>~�_To�� ic��v��S�>{S�%�m1�@lWv= ZQ�F�GHxH{�%��9=]��ߎ�Y㧃�j���J�f�*8�	���k%����ˉ����T����U��2'�H0;7y!�a)i���$��2�z��V�:�g���Q�0��=A�b��;��d;3ih��JG/�?�����#]2#`a��o��|kH0�J�c�A�o:��{��%Z<���
����樠)UYHY��?eS����`c�o����H�`���ƍܒ۰F���7�G���y�_ G~��|@�ٍ�Ѻ�a��qOW�y��)}��͒�� R���Y����w��?V�Ζ�K���|����~;\I����"��k_`}������h�n�r�Ho4�ϻ~|!ߌs�)n[<�8�n��/�~�Ő:���y��t$1 �/���8W�8R��T�,=������&�[��,j�ÆZ�j$e^�NcVov��z4v�d᭫���ۣ;q�ξ�U;����jw/����+![#Տ�>��Z�a�x_��:��㩤Ky|*u�M0�=�7_�J����-ߞ�b�`��o�e2bW�X��Z�{�g���eSnM�-H��Y�����-+���$��.�S]��-�1��+��R���Jy������W�S�*�?3T�QF��
Ї␢�����pxq�ι>���;4n��%w�?�|˂��㾥�iB!�`�C���_���ُ���[���Vh[��t�:'(Œ�՗�Ư��XEh��D��h+���[���r;��F�6а������BcC�闛9d����@�m-��m[p����s���^,u�x�Ӕ/�x��u�NxԞ&�G����������]p�=�B+�N�u�M�ڴYodR�ʡ��䐍�O:fP�6��yU�4����C�	ޗ	Qpȅ�,fD�N��������l1��p�}{�°4�`S)8�P�	�"=A�2�;�����e�`�j�O���=��/��އ�mf��K���U_g�j�s�x�ʐ��uZu����r��=�i�c�$��u�j1�'�m<\��zG����3w�RY��П��8м����r)� `��`�;�'g�YM��sX����2�Amsk��&┑RVXRun��ŵ�|�0I2*���Y� F��y�.#��&��A�eFj'��7)0o�=\X�鋙
�OR�]R5�����(����v�O���Sm$ft�QlIh}fpA��ݚo}��D�Z7�^A#9��(�p�f�YwO���dnդ��c��jb��끭b������D:dNX��V.�P�15��GQ��e~lT�Xc+��Q�q��/5/���}��ǟH��$�_C}��tyD$� ���+͞�/Jj����弙��d�lg��̹
�T�~�1z'V�Jk����]���2�P����=b�R�x��z��'�4
gfS\��b�í�@����7�ڐ��d�� *~�T����hq�S�x�/F����Q��d�l�N	a�r���nQ#,�P��"3[ȟ�`Ќ��g�B��gy=�l�՟�Tn�`��-�r�+����ي�����n���(oE�3�8�6ȋ`˳ b��3�t��K�Y[!�X�N�͉�O�k���j:�[�-�K2+1��ZXB�b8fȂ{�$G�&+B+I��1G^PyVGr.�T=D��uO��7ו�

����Ϡ ��2\A[YKTm�%����'c�!I/���C��y9N���6 �3"��W[�6���پ,0=hvnɠ_�K�h�5��WWQ�Tg +��c3噅�lq��/z�0��7��v�(�_4��1��;M�?�޿��J��f��`���ac��;H��(��#�@���@E�ۺ薚�Ŧ��̪c0�D�u8B����دxeN����F�ǐ�&Jl�O�b1�Z�[�l�Rk��(��Y�Y��͡$��K�Mo��}�L�G���N�����td��M=;���U���m^���La���q���^��b:��+T~yRP��i�= Z��]��Z��Ǯ�:����ǅ�Khf����ɨ׎�;F:���$ЃX��C㨦�������J��޹�6$�2|2! S�d�U/��o	>(:���$+r� 5i��H��d�'�2��>s�`��A����I�R�Faþ;5����@�af�6S�I�)�݌�e�ě�����A��w�?-8f�}cWH|h���}�z�2��G�o��Gqґ6���c�[�62��5����p�DW�N ;>���+�t���R�q�M�;խ}�S���8+q�	L��ΨC�F(%VÍ�b6�k��E��/��Oȵ�p����;)u��{b��m��X����0/`��
C�x�z2�0��d!�^��^�Uo�����|�K��D�k����}.���T�������3�+.�r��h�O��n͋�
��G��f�f��g�i�yo���A��*C-�#bk�\�Ā���Q�v�Ci;"aI=8|�A�X�˘����P�|�w�R9N�lK��eϓ$�O����6�U5�^��z�| >���(���: uF\�Op�����^��,<��d��X?��d&�4N�u�~�EJy!�M��\q��e@�*��U|U���6��vVw|>�n�܏�ej��?^{2���:�������i�Wk/����%�a�d���[�iH/�R�T�q��T�gԶe����	�`Њ��)������Ep!��&-��ĮIٯFT<��Sf��#����D�K�N�0lI�|~�n7��2�G��B\���n��8�������&���3�w���[F�?G����Q��AfzI�@��J3kO41�ݪ���'����=nMń�{�j�ڣ(���UbF����J�0�X5��C�x�:d#H>�$�V�jW�
��N�ӱ��6֊E�;0�Vˋ���JK$�,#J�0�P��ʺI�{�C�1�Gu�VF.@B�����Vd�[�@�	<���8��P;��D9R,$N�+`�������H��c�e�jIv���#��Ӆ��Srꡧ��$��*ƚ)������  ���x>��Ȳ�B}В����_�a9R
��	zI�⋩}�2�����c$Κ�6���Z��k3E��M�[j���` �jT��� ��ǎ%}��T<��5��1^H���B��e��t�
ɽbv,`�q�D/���&��<J��e�C< ��s�k�6�&�2WN$���b�z.�toX���O0iIv�� �rࠢ>ӓ���ˌ�*h㮝�&
��B��#J��WMv�I���bcێnJ��t���owe�+ �n��ĭ�fu�f�}�ӟ�n���Ϫ��ee���c���N��+����B���B��2�EK!��[�H#��x�)�.%�����ȕ��m1�F�ŁCS�.,Q���̾��*����o���)�t_�l��hO_��9���3��}�KP3��]����B/M�S��A�*	�ܗ�C(��E���68��*���R4����E��W���	~��P�F�2ۼhE������Hz�Gtsӏ0��ad��:���GD�V�@��-�tOV�<���s�����~$�p@+U|��.��8#��ԁ����c��+W��y�V�6�Kp�>-�lK���g�`���\�����V��4^�	 R9�o�r'}��{�l�>*������J��h��V(�O6.[`���Q�*�eIr	2,I���m��^�T�t�͢�p�,��$p(s�:XNL��zU�WS��%�i3�ǼS;�)�$O=l-�&d��X�i[~c�d*4����8ڂ6�.�N&� @�͵����%�-.\�0X�t��|�ա� ��x{�ݪFU�w�j,������R������/�~]/a�@4�&L�!8����+�x���{;��� ���=�7��6cx�\�("� ��oKz[8����2!�us�4ב��`��y&yh�~*���m�#e�[D����EYjcv�-1��#;������i�K�:���!��7�da�ꤝ$6}�v�|��e�7�L��]�QtP�X�]�2f[��a�}R6M��}�2gc��JQa�B����2��������s!l�Ռs��=��\N�j��3�d�Y���rͧ���m�T�b����S����j&{u��'U�(��5�sS��=��١siQx��S���S���U�0��yo£b��OR4p/��ɼ�"<4�� ��������Oe��%��8���,�3ﷱ���Tvx�Ib�:�}t��H)o �/@����ȝ �ȇ��Ų���.�R �f8��|���阔",�/=�:��#�׀!}!	o�n-)ɾ/��3�Ѷ#l.�A|&�nǆ1v|i}f6�:+����;��w�:f,+O4�ٰ*�����@�l�J��Paߢ�#�XT*��j.Jh%D�eS��C`o;�}�Rxh_B02�~*U�9��yo�g����	��
�?��0e�-�-���d����i��u1]w? �([�:$3����a��!��B��a�7��,}����"��ġ�=�m��q|0��"�ĳz���V����c8m�=�-�&"O^�־S�����ʭ2v.W@�C��"^W4;1�KĈ�Z�иm��@Y�V�V.(胲K�AM�:�;0쨇;��{;���7�A��7�E�-/�)�g�U>u&|���%�M50f	_KJ�S-[��� ]kqu0������I�lb����x^
z�HV�r��}8;Xޮ�n�}S3X��v�PĄ��&<�ҿ�A`�8��;�[��y+��<��
�:=�"�E��R��}4;�h���=�����o@[��5�? �PT�E�����C6L��o2��L�.b��_���Y֔�$�*�Si�K����eƟ����u��"�+��<�:�Y#[ޤ���k��&h3��>��l��v)�b֪���a�K��q4�i1���+"O� �@��`�?�p�����1�l=���D�?�Ш���
����项q�J�B��L���@�\�`��;!Yahq�'�P�]e%�)xqF�{lc���u�O��ft;}�с���1`"O�3}u�,yO��]�OW���4�f��yR:�:�b��hu���Hc��(/��(N��G�N
��
ˋ�~�.��8�%Fk���=����-
�T����18����f�SHK����d�
I���ƪ�3G\>~bkΣۄ���>��Xb�	D��܎�&�	��<�0��Y3�3lu$��<_@"Qj�s-��h!����l.6!�������v�'��d���3��B�(8[^^&��͋�?Q��K�+��Z��mD#��)F��=覾���[:�Y"�<���^�q��^��S��Sx�ު��坦762�_A����~�]XnVl�VuD�w��x�5V��>���Q2���Q�p����a�Gfv��Gײt �t!dAX#+l��$#�rHI��k�B�5m`��:�-
<����z��8�� t�����^-���smp�,��W�{��jf��(�t�ڪO�­�DWyR){Ιh��r�O)(� a�%Y�<�}ᚋ���)~$�����$Kv/�%����6�շ����[T�~��U����6q}�O�^�_�ƕ�n��啙Q�$�8��m={�/.���5�^Qdv�w�����P#K���Qyp������H'@w�oE
�VM��G���x��L��B��764��g��K�� �N��UJ��&�V��{4�b���ٍ�}ܓ��"��P�Z�^c=�w5k�{�^G�����.x��k�e
��G �J�B�!��0�[��}2B��=��Q|1���ƴfs��XfİB� pX}�Hq�����Ƌ���r{p��n�m,��Uǜ�v�_��MP����4�����l�������DZi�����o�7�_WGl���`��zW���]}�.���~EWC��2D`��"�1*�7��>�F��$R�h�<��(�w#U����%ǳ�WY��`b_Ӟ�^e�G&��/�6����@Ң�mXK�e�&�y�d�0��A�4�uu��~ȷ&�����U�df�X��|��>�}[rs�^�j����7v�>9���l��չ6��@��������M�NPL�ز�|���)H� "M4���W��E8�P��pc	փ�M���4�"�m	�I�����9ǫ�)�ŝY���������Z��`�!v��p�&PQ�#RA�kn�C�R�Bʟ����Q;�3��V����,��E��*�HQ�X^=A�U=���DvZ?0��m�9X2���.��Z�ѪV+0�ٵ@ۼ�FϤ�t ����!�%���Lb��*j&0j6��$9�� `m'>yR$�Ӡ�1"�?��F�b��)�ॣ�:uU�S��Y�����wN��2l#�������n)5�B2n��,q���z_�����,�W��op��n֡Q+�ŞsF�$Ӎ���}�!�ձ���Ĝ�'����}��BxP�5J�@�KѴq>w���?��9���`�7z�o�:�t �m��&�Z��Kl~���״�	�]��nڶ����Huڱ{M2���a�W���K(���R�^6���ČUPK~FX�?
)M���\h�����bX�G��h#}�B����t��^���w(�
.�X�t����-6
WW���!���`6!y��⹒y(�ꢈ%JUu�T�c�晌���<��P]��C�I��I���KQwJ��:0�b��w�;5����W�X��&ﲟu�ӣ��	_Q�/���-dr��o/J�`L����LM�E�W�xڬC��#��̚��Z�(�a%A�nI�[���{CK76k��Fk<�I'*�v�=��0��Z�&�W��f���貤t���E��K�VI~mؠ�6�3� ��X�4���Dicy����(ͯ�b�LmO�X�o�C03�s�f
2������s�"��>E��{ϰne�h�s�����w.c�n�?N|Iw#tP�NY�*s���7�Y�~�|�:j?�vB���(J!��b'm.��xb�M|>4<�]��x�z���=;�~�-M�@vIJaUfs����?�)&�jK@%�4��X�QR���f�������ݞ *����צ�4��~����<Sq��:渠D&F��������� C�2������g�Y�5݂��/�o�&l40ce>	Ќ�C��:�㉉��JiE���Z~�
j�5�*Q�a \�:y�$�DXcș���"�ŕkb\&�<T��0_S-�����zt2����[��yz���%��A�<v'q9��@h�d$;����E���b�H�u�A�|_���a��Q��Q�|t�z-�F2O,u=�.�N�+؛1�3�;��(���Ʒj=��w�r�l멻wJ^�Р����9�t6@�H����w�3�$n.4��wK۬s�?�:<�cr5x��c�濑�r�50>�x�f�2��i"�������dQ�Ǫ�s���L��S�k7su�T�{1����;�"�~����R%
���js^B��c,��g��f?�)iVT����q� rO���B(GR�]��ſ ��~�v���n�&�X���HO��A�F��������ط�����FR-|7�ذ��F�}?_��~�c����U���ݨ�	4���u���T)��m���_Dt9�;d��P2�T �_$˭�ئO�`M�^4.��`,�ތ�""<�Ȗ��H�Gf���2g/�L
��Q�Q�+��9j��i�^��D��0_�B�D������*Ox���yn㊗� �7*�P�K����3�U�>V9���	����M7�j��'�zeW�|�f���c��D[ވ��F�&�o'9pҍ�H�9:2@*��h'�)�Hy�4��9#���$���_�`W� ���@p����ኹ��n�K�8,�tX���_^�|�K�q�u(�߶I�U����,IW���a�	ZY�ݘɈc��P`u��{��w�����!��Kڨ�<��I� ~qAw:��~���.�09�)y�*��z�p*e/f=o�sR��*��mxi֤i���IMOLx���'Բ�[j�a�
)��&�2ua�ʪ�]>56�O�IA1�,��؄�k��v��"RZ�@e@LV3�Aje�i�L�d��?��lB���3J�����?\�;
~�)�&�V׏������d
���\e ���0��[�$	���¹�k挚x��"Z3��0�-��b{E:��d�9rj�v��縑]	���6�U����}�ܘ4�cQ�^�0m��[�3�%��Eg��R���}OjG���)A�?��)"�(K2H(�CA^f!xb���S"�w=	㶆��JJ�+�=7Y�V�N<��Wt���I�aYּ �~��d���v��q{3د��ơ!n��R�G�+8�>�����!�Ƈ�,_��snt�t*���؇�� ���ЫG�o49�o!�cyN�F�V��8�I��ך�{1H��Ll�5��kq8
\t��m݁���9z ���%��#��g�y�p~�G�<Om.��}YQ����7r)���!<0��}�C`��t��Y��"#F�� �W[���"��fZ��=������&&�c��
�F����AP�pN���q��J�9&�_!g��k�Mv��p�����b.�j� �m=�d+���%�y�������FOW1*Z�Ɲ*�I48�LS�?�F��y��RY�İi˾t��ħ��Lb�u�����p���h�3\����o�o��[�̷��T��3+Sp��8�ߜH+��~xUJƨE8�NrF�v^滯#e�0	�϶�j�)t��a����p��N۳��%2{K��V&�f�2�#\��eSx d��OUP��]�uJ\�W��&'3����D�a�kx�3��Q�Wzd?����cS% :�R�/��l�f���zZ�RAxz�z���H�e�j"��c�)/��ޟ�H �݁���2fwJ��z��E��s�����es����Զ�_E7pI�Ъ�=���h55�;uė�n��X !���:�c(�5���q6���G��8[�1��R�9�&?C�ev擓����{�
xd�}��6~�쑭a�g\~}A�ט^R�������+8v�:jm�^\�g�Š�G��0�o����>O��p�v E,�N�h�=��ܤb�T�$��
>0b�ğ��<H9n�����z,�<�W��|�b��c���Ȣ%����P<?i��Y+���	�m�%eC�鋓��lٗ��{�����]���ݨ7&��O-�Nn�Uz����i7�l�n�R�����u;�x=��vq12C�3�6�i|xKE�b�f��e$!���T�>�%�E%� ���'Q��!=~����٦����/Ǆ|y��ѠX��̟T�8�5���;o���3i���B�P� R�[{��2��n�~�_9�8|*y�e��>����J�v��;��'�rs�(ì��n1Z��gn1,⦮F/x5�^���/Dp'�90�&8q��m>Þ���L������q�8d�!����F�!��]�#~(2?3 ptJD)�Z+_�(���35��Om�I���ˁ�<��� �kn�b��O~�c�-JݪF����B�:v�$�\9i@"4\A�p4�yu��FHEb����D���B��#�*�u����8Ǧȗ`aQ��>E�7�=���E�</��c@a�� �^��&��o�3'�ׯ�Z�1��jl����d��ՙX�~b�S�a��џ�E!�V�}���ݾD�l����SF	�bȯ����[,�a�*��j��[3P�@ռTO��F�a�Hm�n��	�Z�����vL"��@�
u�ސ3t�6�!�d\������Ըh%NR���&E�"i�3��v+�
E��"����.�o��1Γ�y�#�6X�f���
U�>��%�ۧ*j#���x۴l�N|�e��M8������/�����/���7F�^A�i�;v��Jz��;/
+rE���vb��	9Q��G���1_.;�[�ZW���P���[�&�N�6��ѥZ��0b�IH\� ���hίǧSvhuN�,�O��g��V��9RHN��wIfʐ�UB/�����[����ir %�mZ0a�b  ���w	�K����E|�<�ڻ�'#��~/���jR���/�E�4���"̋�4XZxX��H@1�G$��6fؒ	�d^t�,���^���)��+ an��<��쵘f�֖�{|�ETlpgyU�#���I
�x�>���F�_i�{��Y����W�L�~`��c'��/*�P$i��0�(ОZ�����@�$�-bc�����NgJ�kTc��p>�1�ʐC$*�6o��Em�5E�mex8��a2�+U_ѕ�8�×^a����x�5��>�5�B�.BY:�@��=A����/��)[�)B���̮�jp<�%j,WT�{�b�߁$�p)ٯ��z6��S~8�a��8`^P��w�̰iD��a:�vK>e.p�4e�y�$K��TFe����L���*��{�Z3kE����Ck̡>n��`B3S�b�1��d�jOy#;-@"���X�A�^�Z�R*��Qq��_�?���+��H�{4��%�9�!{(�똩����������\���#��B�%�ڶ��|)���v%61�x�Z|m���S0GQ����؏i����O�w��P�)�Qp��]��<Clw���p��!7��t���O��8E|��c��2��a�Ŧ�����[�i�R�>�ȸ�������òfᆾ���$A�/c64f~�V�����C+�u��}H`Kc��ZL���DdUŁ�}1�=f�A�^6y�������o��b��a�0W����o!E�� s�4KBl�+A���.Wa5����o8�.����I�L�ؖ�YX��/��ᛌͿ��9*q���W9��hE��N�_��Y�Y�4ƅ�J��/.�=Ɔu4����`p,)�ҠJ��B�1����G#�� ���tOdr��*�6;GUDڎ���6��/�?�bٶ��W�gdA�^�����|����ipўm(KSj	��N��ذE=�ޢk�^`~���B��+0LɊ�%�RөX�EG_�U��y�Z�|��X�*��!1ujH�
>�9�Aa^�-�I��œc�>��R�r��(�[FX���T-V���@�IT1��Սh��PO�{��O���Łu?���E�1սØ�$b�'ݰc�^7x3��nƾ�ծ�U)ќ��-i����h�">ׯĄ˔�L�l��0o"��3�z�"�p�Y|qaA1�gr���,Q�ט����v4�ɰ`���] �uy�(�O�gYGǤ����? ܃4�V��a���?w�J_�~/Y�=��0���lD�wP��Z�u�V=d���y;l�N�ZsӤSx%��U�P������+D��g�Cn�=� �t��zQ�Ls_.�T����'��Ϲ��T��QǪ��GY��&|ޫ)�3�l�|�َ:p� �����B\f����bٯ����_�8۪L��d	W����7���Х�b0"-ʼd�D���&�����+�7�\�$�OR~{��ř��� v<^�3�q4L;6�
��9�*�v.�Ii��%��!l���?� ��'䌊�YK�9[<o��R)��@��2�����LX8{z��./�l-��*�!������玒��,{/s	�C2y7�d�J<Ͻ]��==`�����{~Y��+;*�3����N��i�D�$E�%��֏|�e���-����5`t������t=��Be09\�&�̶���\D�V�"	S�ׯ�u��������S:�����g�q�������/�a�>i0�Q}�,Sާ���B�h =`S��hG7>�FY�uI�A �GO��R/
�acR��S�g�(cTq�`����7�EӋ�g5�-Z��Z'0i)�c�?	�Ħ�ɭ<�G��Kd�����v6XJo��I�(]�bOnbWv}kF��R�0H7�lG>m��������8�i���8/F�K��O�=�������%�.��M�SW ]\��d�)��LK+����%��չ������X �z�t�e�d�Շj=w��1~�4��8<��w6^�p��ҵy��,u?4(�K�2�q���	�u%r71�;���z
L~�Dn�Ԑ��R����5خڂ�ˋ�̆�<nr�����?��
l�t�n�ο����NFD����a��ɲb��otg�M]�[uj���>�L������k!�v ���шj8���M���M@�ͼe�&/L�OS�+%�t�������._��
ᱛ@@r&Y7�o�%YF˔�#
��F�z�(,���Y� 	FI���.'�Q� i]�w�0�q�F�3�e����7��e�S�Z��#�ʢK��q�7��(�l�Ό����C�']���E�/��ₗTO��盔�m@�T�/����I+�s�l�m�7X�#2y��%r��QM��ހ�-�4BX����j�����@|�S�G1\B�@���� �^E
�N6��9����ەx�A�?F�J���e��D�8!;��jp1)^�.��Gٯ݀5�͋��;[�C�{���s��N�U�zy�����R+n��$�����n$��@A�3 /YQфXs��`�9%�ǫ��~!���g���EhJ�߉�Ú�)f�P�."�Ǖe���WMT����ׇ�P)��7}�PӞv�o���mZa�q�O 8	l�c.���G @�QmрrA���!JT����(�#Q�&u�c��L�)1��B�Ր��S��5� 	��a�Ѐ��Q[�h�w���(#����gQ�Z�������4x��"�v��Z�2���&�lyt��Ꚇo��(7#�F�qj;�� ��������m�$��G)q)Qm	��y��K�+x��P�=�CO���)76D��È��?���ED �R[��pĶ5�܈w'�.�����qpU]i�F����{W�$%�L��$�i����Te"���?z�F!A�eW'����{��_���%G;[-H��7Jpj3��d<˵e�@YJ�d��Z\V]�KDہ"S��~⬙�yh�R|ט��5�X1����� �P�)��%�(UF���?yk�T���@h�86`P]��WNL/`l1�챹���7^t+
��U�p.y���hq"��Zĥ.�=��t����:��XC��㮡#p:w���
7�G�n[�('x8gd����YT�>S�b�e��Ǵ�	�X�+	�f��:՜@:�]9�w���R嵠٬�l�>'�}����VTפ_)���)��w��k�0��	�~W(�Q5O���_��Rq��L(y��{[�Ōw�S��m���q���!�P��K�U)���Lإ��+$��R��3h��3P���-I��"9Tj?��,��ԋ��ѡc�"RA��H����=�kk�ɘO�+�\Ľ��S]q]���d���X��[|J�X<|��$,����cl�����\n�=�XAS���Sxݨ$�&��K��L�/�䙃A�5�0�v�Gk��e��i����| �����
��Ƚ�V�lO�{@�
8���e���e[��0pd*%s�CS)�O>s��R���h˧�Mݺ�G�b�	�7S�I�n�������0h��-9O!5�����ק�8����x;Z�ss̔�!�/�rG�Yz�z�\�	�` �	�Mě�Y�Wg�o��Ȓ���@�Q�[�a,7]�qk׮P��Q�a��.���*��i\�>���}l����n�a�Ui�Lᚴv~�'So�w�Gh2��#�z�Ʉn"+#�~Ԭ�S���mW�U���T!��ف�I+�`�:���|�-l~�e���|�p�`0�������b�q�hL�����$u���Ȱ��(�C�`N�e=|��$J� �N��(`�M={8�3륟8{z�8Js>3o<����O�������X9մ"��i �H�B	��A�n�(�:_����\M�[���G:����[7�b�Qh��q^���^��V�$c�g,IjѬ>\L��~�j�nZqR�F��R�_ܬ�?�xV��'@��PG*�ޕa$�~`;��V�4������/͖0va��@�pjl]����/�e�¯���US���C��-��ݍ�?&c���^	[����H�q���<�%�g1јdᏎ>,���΄�h�l�j$���I�e�2����{��a���>����N�ˌ|t�t�1z������q�`5`�`��\���9Lz��-#0�2"4��J3�(ejyۄ�b��D�Q���:$K"�vA��h�z��<NH>��?�K�nt��Hz_j�i̎��<",2+k��0��C�&
�BS�)����jsa��Cz�:����r+5 5�xlD��l���n�6ko���l�n�GKG�xt% ��=N��2~�*��/D�[#�Oc.�@���/S��y $M�1KW#��n]�T�s0l�R�-𵜿�{����<���E2�rh9~��eVz��%��5?��6�/�,Aނ��� ��Q���vJ��i��C�����QI ܢ"�B1��Yo�R���}��Otl�;1�F��XG1Y�;j�=x�"i�u�W�]!4t�#�4��D��HqAU6=x�<��;�k廞W	I�B}�h�m���J�$�����B���� �׏���qzX�������t]�}tŨ����o	y��6��. k+b��U����X���.���W ��L.�y|�p�%�r�7��#S<9���-E�<�>~�� �����1��62���W�-fn-��q&l��r����w�p�A�P��0��xR"&NWR@��[�/�J�A�zx/���*��p�+Pe�%�sns��n�H���6���	�V�xD��=#xez˓S�[���g.˟n;c���r:$�{�iJ+�Tn˕2N*w�=�������2ˣ8���]�%Pdޗp�)y�M�֡�����]�E5k��\Y�
G%&a�)��*�uԡ�.!E��E���6l��pv�&��I[��!O�v��@�a
�=�6w�$n��Ӿys�*���=��#'��m��&CBB�?�I}����w��M�Q��j`B&�l��s�
�1�W�7n��9@����Q�'s���^!�U�+e�+^�Em��D��{S��=�[�h�t`�\J�m�_QV�	\��KI�C<�Ӑ�R����V~�#y���N:�ïգ߀��K�3V]�J�XN����w_���>u����/�u���Y��ts\؟�<Oנ�r��d8��>j���UA�����f)��n��Gš��)+?����ěD�D��� ��h��-v�P�ı�;�p�!jX��t(�ښ#�㖑O�#楔<���m��zcM�e�+/�l2S �5��N����Npx���N�X,ͧ�Y�ʐ�]x��t\���ݍ���h��_��̃@]�[W[Qr@�	&�lM�}@�#(L>ͭ��E����h���o�|ogx�4����>���~��4���p>3o�9�pضY��^��S�ϵ�"�_���u,��0�U�4��\0��pP'��iS��o��֎
��EA ��g�M�J���W�8�������"T���	�5`�4�9?��� O��"G	K�S)�:+4E=��1v\�l��u���4HSu7�xS�J;�(K�5/���Ɛg����6���&qmca��La�Q ��X#��3k;�z����Kҳ��=��C7���`$�ڌ'�0�O��!	�^�ygR6�?��ꎴ7"iz!oyv��hK!�m�T�=�4Q�ן�ؐP�b~>ϝ~7���2�*U!4s��# ;�U�g4D�#�L#7;XU��%{�.U'���D
�������C�	��=���m��z�na����.bw���b
[q;f ��>�C�ǹ��Y�]b��Y���v-e���籷f�C�+Ģ&aiӍ�:��)j��0@%8'��Z:?�*d��Q��m!ɑ�Δtu����� ���6��l����C#i�(c�S�;�Pt�I#[�KW=j�}M= ���B���,{(�fR'ٞ�߁��E��c��Y8��dg$AU�w8�p��!�Y���=Q��Z���ú�:���gM>"pA�XS�q���c���c�w����a��������q%���| 0�����5Q|��$\�m�MwB�Զ]��P �B�0����#��M��1���3�b�寧��>l���*���ia�F�
��$r$��8A
y��� �FGD�|��HB�P堐P*'3tX���e�8�����H�<E�5Y�Q�l{aw�<�����b�~�I��8����f�������$�:��a�m�N��\ܷ9�3 ��2�[�r�MM6L�@�wK�?#{f�[p+*Q;��Po��p���V�؝�{΢"|Y�$䣿[�Ņ�6wZǧ�Zܤ�H^�, U�A�Բ}|����}�_�2�=�[�wă�SGp�����#��O��(`稺�&���O +�3�F�3��]�.0ۉP	a{�@<BV�!��Y:&��T��ʂ�����ְAh$-�=t�����4� �	no�4����]�:��//Ox�X.Ɩ���N�"��ʽ��tC��h�grv�&���i�� Р>�.+�!��Q��h��ϰ�����D�߈ai�U�I�l�������.���A���9>�i�Q�0�e�;j�QOd��%���٪~���U�\ЭFE�qCj>=)��[�6����[�׬0a����0z=���j�o�$0�,<�nA������8u�^2���%��V?3�&�*0}�f�np��/�{*`�+�$�����@�H[K�^��z�U v@���.��N�Ǣ�$v�zۋ����a��WZ�h��M˹J3�䚨��"$a4;Ęo�
uMQTS��K������i��;Y��_\P�y�M�S�&�+ׁ������dK���O�����dj��:Ϥ�˽R����y�Ni�  ��3��s�*c�+�ZvVD�]���K������G�*�����2��S<�t�]��Xf�Q {�nM����0Q�p��x�8�'�MH�}	��MEkD'B�^>�Z��&�*.������M�H�R��H�\LK�Y�Nf���5�xl��rq�����2|��Z��*�YY�/�1�3���M�ZUy�֤���e�c��~�6�[������I��u<QqL�.��@D��du�����/s:����yT�\A�d�uc��ſ4�NV�ZBg�u�{,N�4�MDm��[��8�K��dL�4d�"w¹lqj��O�[b�Ui�䃻�_��
Q_���t
�w�ޫ�&,��yd{p"�>�wJ�e
��Ϳ��i*�	Z�ϲ��a��Xؑ���c��܆ܧ��I�hЁH�d�! |�0>�*�jWl����kn4��P����%�@�(=���r1w<��*/hYĿk��w{����S)9�-E���fJ��0{�O�MW;��d��0����Y4��AZ�6�^�����oR��z6i�wH猸����5婻�S&��k*�C�ȋ����nG�B_(	���cz^���v��#��JW�~�g$Z���2�L1�O�а�!�c��z%;6�r0��"\`ԯN�������F��Њ}aMA�	;�N���%�`���\|K�[N�/�q���Yo�(s8�	��Ӟ�"��$lSpQ�u����j�'���iS^�er�v�x�-������u!M*W�}�F��=������ޑ�\W@0��PO�YK�޺��s�w\�.ʹ��
����כ�8����q.T.�w0��*��bXۻ�m�Ǥ���	Ё5?�`F�Q⺀�k�SgKo��;���`��I�	��x��c��(�M=��#�lX����<���y�z-MG�^�hA���Ic{���|lp��H���F�W,4�^���yY����7\�U{E��oS��M�ق(��u�X���R����p"&���卧lu��c��c���2���|����I6�k(UЧ����[,Yqދ�48�Hc�=F����lyν�_-'��Ёv`�y��b� �$"I`��6j�>wC��D���\�4��6ݶ��B;X�?�)��G�>�%ǐv��
��xtM�@�5�\����)�hS�B8A�G/��/n��33�!ٴ��nr��m�]��e�J�/����Ӂ҉����c6$�	#��5���M�_�g�(���Kl�Lv�n�ð�1�X8s��"�oN��pwA��Q	��H�v n�����C)�#Uq�b`ߚ���rsMq(g�x�v�Kȸ(ᠢ^4>5�a�`�h;�n��}�,+�y	���rN� ?K�)1�v�:�!}�d�T�o��hy�f�=� ϡY0�!�OXQ��>���ɑ%�a��{�����ʺJp�$��M6�Man�-� ����A�07!tg��-�t�8K`4V^�s=ρ}�P�/.7w�Ϸ�9���/&�#q2fߟ�k��?�|�֣~Q�N�4�6��HC��(����ȷ�%��w/��b�����(�@�m�����jPu4�uF0�����^?C}/V���/v��TOI� �h�����uاa~+P�v`�k5D��Q]	-���櫭Len]R�p�i� �O��y�)/uj}�Es��ud�4�>rAz�C��\�א�%N�.ډ^�k�AE&2���ED���!��W�y�+���^�v��]�9o��{� ��-�}�߂�j���M� �o�t�bpV������!=���d�7�ui�ͺ�v�⺘�֪̲#�s{�n����r��ː �7�Y�ߡe�{��xS�:&�,VΖ���i�"a��9�9Ze�L���V"�iR��܅��,�z�� ��8���V�d��ÇT�`�������[E#a*��͌yq5�/&.�E��8�X$�H��Eڡ�$�%|%�i���h�G&��yb+�1�{���f����cc�}��0l)!�L����@��fU�����>r�#�'I� ]�b!b��w45�dk�8"
��8��C��lCRq�,w��C��S 8Fj8�^7��k�ɳ�p�Z,E����[�@`,��\mF�h�_H���6��6%��S���k�6��s�A����%�UvoɁ�ԝ��FGQ�lgu^6(�3�h�e���cj���D�c)ǀ�~�k�LV����6i��4!�	 &�1D�e��-M0ì��\]=S`�kC�0<��J��ut_�<�M��� v�p��
ي-׿�r�9�E�{%����7��YM��m�y"Q����,��)�ã
�+G� r!�V�����o�eR�j~o2_��N�`��E�~~�m�d�Gζ�)��!����x�"s=Aor�@l�@:�D��M[K~��e:��~�_�k�YW�����qY<��BQ�~&<��S�����ȶ�]�E�T"���Ip���%�$8�X�qyZ*�u��Z����㉣�B{ϼ��d�n�ț��e�`�G=�Kڝ�$ݷ2�9=��h�%���}[W��	L~(N��
�` �S��Y��N��~&A�ܚepoy]>z���48�)C��K�)j>�W�*zɶL��U~�t����*>��s��g��>�!~#��;{�����>���/ٞd��f%���z �)�%3�9�+ib	�3�����0 v����jӁ,������q�:��M���Չ���h��󌢱�<1�3����?(l|�?����Co��9:PH����
�e���{\9??�3�W�f��K����逿�Z�i�j�ʝ�����e5���%�B������7��P�S:9ҹ�5�e���"���Ϯ\
��ɔ"�Q���mv���n��k+�� �,�G��
� i\����b.�V�plgqY�u�NY���WP���\�)����}������fz$�I�F^�w����?��s&�x�W_���`���5*�E��H�9K9�s��R�M����ߓo���\M�O�bT���S0}(��j=��mNM��	��_���m3�_����#�Q�/�R7�p��oŞX"�����G��P��pX�#4�����%m�g��{KBD3����t�:ףS��Y�c����%Es]7��)��������E<}����՘���m�nNI;�D[��l���SB�:��NH��s�K�	�Z(ܔ�Ȳ<z˺%Hjx��:9��֡���1ڱ��4�h��hg(2���I��F��ff�Y=@��Y�$'G�l@�a���`�-�単*�D#���djdզ�[����ٚ���hzlMr���y��b������:)Ղ��q��l�)&�LwY��CI�]-�lB�X��˷{������	f؇�Q��!�d� L�5H�F��Lg6�yD��a^�\��D��X��K��[M���"I�){F�Σki\xDs�7�_M%o*U�16�l�>���|M��_f�-��<Y�*�f�un�m)x�TsZ� �]V���!�Z�)������� �͕F(9J�C�:���V��������I{�C�X�0����ܨ{g&ߵ,-���:��a���XW���pֶJ��G��ޫDZ�->U�9�~�����S���B����d�b^��L��[`jAe2�Q��'�]�.ߊ&2�D0I����Y4�j���,BN��A��T�Ά�?ZZaK֤Wȋ,,� �-;��t�� $�%���fV����:rHI�j��D�[t�����׌��gC塽��gr�肣OfR �b�&˻�)�h�l*�v�_\L��%�>�H������ݰw4��ʽ+�eA��_xဃ��ta�#��a����jA�/�÷�T��*L\)���F�]S�U �N������O�z8�S1R�-d7�X�w$ì�Z_��B�*f�<KR���/&d�]��:-�p�Y�I�����g�qN!'��1���0����mv��\&
��h�M�e�k-Qx!l�9��1osԢ}A��Y">��s k�L8�Th	���ƙ5nl)�1A�"g����HQn��ٔ1W��Ys(��h�R�$sdr��ϵ݋By�'up���H��Pl��ו~
%M�L���AӴ׽g?�D�}�ϼ8��Wl,�����@��	@F�#�p�V��Ҹ�Ź���(-��[����j���r�?���Q��tp��u>����l?���@�S0�@���,JpP�i'r�Ȫ5���mA�lpur�B��T�r� YShsz��Y4���F�X���Ȝ3k�u�/���Շ���S�	U-S�5��~��3&���f2�S�+�ڟ	P��>Pݽ�S���?�Ȕ6��O.����'��0	��X|�W~�'����FhG�;<`Spbp�m��/,��Q��C�>a3m>N�/����� ������e������0�'�C҆V&��[�zB��͌�ER�
U�9�@�~��#�����)L$������Un@!�+PO1�Bc��@�(x�}0�j�ݣt�:e�9�&o���?C����D-�/��� �!�{Ff�!"�g�O&R��YJ��*b���T�_ N��}�;��ܠ��&�4R>q�ό��,x����q����K7��j�Q�2�j6*�����ec"̸9g��j��%�+ ���%#�����gGG�D�	�4�?�q���'�D�Vr�x4�IOf����e��*~�DB��i*RY�o3�� D�C�|)�����2���of^�vm-a=@{�D0�E�5��E�K=��M?ο�+��O�\�;�R�s�b�&r��{N��M5Ä�	V~/7X���vֽ����}�%��~X�︖���pCC!�J]�,}DQ���	�������ͤ7ɀ&*F[���fON�Yy��K�n�.�E���sv{^�Ȟ��s���L�ճ?ƨ�:j�?�e�]�D��::I����K����U�t�t/W+����휟k��B`	zñ#�Owܦ$�����06��ᒹ��g���+�J���%�\Ӡ��6�IR�8g�@V�n�ǂI���s,R*�W'Mod�AA�c�9} lT�G�����:?�E���?V�R��� :�pB8�������b��Y�j�*^��9-��Y겮W{$����pu����6��%'�ڐ��s��I��$���Bq�Ft�2_��vh�{��L��9��O��oɆ��0���j�3���G�!5����Y&l�˛x��h���"��o=������מ�t�!m��}��H�(����>5c����\`s~�Ũ<�T��F��p�ʩc�u���wQ<���l����fX8�Fv(I���&�i{*A��q�N��h�{�)M��" ��|ޡ�@����Z����*�pf���tT8��Ð(%���U�� [Y��D��wW�
ɏ���|��x8ѫ74mh����jx�懾@���Cn��������	�trq�J�r�16��{^WI�����}�����ܹ!>:ėxC5d�o�&�7w�l䷷�
�9������,�#���y�#�dr�1��rk/Y����W�S��
/q
�OZ3�!W��:�xOYk�VAQ����l��Bp���`N^��K���_�C��P���8��kp����f��()i,s��ːv�m�'PB���9��P|̜ܳ��7$I 9"m���P>��4\m
z�&�6;���bV��3�������<-Q4��@�.=TXv^%��DS�\6s�H<zQ��X�
�?P|ǃݼ��(�S'\7$��Ѽa�A��ŭz��~�1L��b�4b��-�_u�l��/X{�A�w�<R�������F��ݝ����L�@Y`%$�P������`�|�����Cr4N��'�>ny�g�;�)<L��D��������az��5���P����%U �=�%ʟv�x�פ"Wt�x{qr���g0���A��w��e�Z�{� ��T��ճ�(�v������5�zL �,(MJl�s1�%�D��j?F�F��B+S��F"zG@fJm���YP,(
�4���Ւ7c��8Y�sЍG��x��G�Kr;���G^�.����V�߬���/�������z�OwO5s�n�oZ/Å\=���E�;�������e�HTe� ��؏
�Z�_Rf7d1J�}�r�o4��PIK45D���%T-λݵM��*����q�+K���>Z�nSq��d	9��KI�/��ߞ��|���*��!����&�4�7ҕ�m�v��F�V�* x;W�\�n�
��8b�.�dK�������͢ˍm$ƱUx��A���_ʳ<W�*�%IN��ṱC�c�o�CS��ɰ�y�d��${�*n�`�T��Աȱ:�t�:
P��ڶt�O+P�q�`�l�7�j1[�v�َ�~=}n��!^���1���7��r�����(:��l��W��o"�+�����p25����T]Omt�e��c8a�ñ��-�.BWO���,�}���p�J?��A�?>�4�!��B����	��r��w~��v�~��BL�g�㕚�����U{v�H_�I�Z�O]fu��!���!@*(�b��KȘ7�t��t�Ю��|��f0��
�#�a�R�K��H����w�"�����AŠ�y:�����l&gBx^C��d-��/�*�jdq��UP����rn�[l���zc{����G�����GFfR�������m����J�ͪ��I���C^�2K���e�j�E��Q�R]O��o���{�urj!���q�r�uő4dJ�gu��Įm$.MA7��vм�X���\���{el�/I! ��i��M��_��R�>������ӹ�ž�4�c�f����o�d�.�b��u�}{"�.�"L����Jx�o��#O(<%���`b�ms ��Р�K`�<^��S�4����0����Tכv�����]EaA��}�qϯ�L�4)��l�Oɡu�w��	|kf�jrWq�~�򬭥��Ҁ����zT����+n�)�>Ώ���z��:��{�{\��|"������|'�i��D˺��y��h*A�ٖ$V�;��
��0��;0�0'�ʝ����rΛ~|dH�;�֪Bz!3��&S�ɝ�V@ٟg_�7)�-	�a������ė6X��6�����a��GOe��^v��5����jπ�U봓�RG�p�_�S����5]�4;��t!r/�H�OF�~�*�lEߌ�c?�QW��M�T�2be���� &���oL *���׷�^�Y�!��������Nl�X����%n�!�^0��L/�(zÊ9�2����O�R-��*�v��niT�'K̼�E�\������\�ErNC�ε���$El
S�v��'@y�
3�Y��Ӳ�9Z/;i:(��X�T��M��)�R�|[�61��
�C-��\�yU�s����T����+%4�ACC�j�'}z���.iऺ&��Ж�3-��v�N����B�P��ޔH��~�پe�`
-ֽ����ߋB$�2����տ bY;`�1��Z,��h���}�"G�ͼg0pਂo��H\���[ ��n��(3�)V^t�z6Pyk*d>�:��/�A���h�Y(�a�w� ��^�~���� �([�L"��tG��"=���dpaKF�ҹ��bi��ؾU�Z��B��[���}�������S���{c���pLZ�3���"_	iD�����1�T�
��sfCX��?Μ�n�pE�����!_M܎Ne����iz�pO���٧����M�>f��s�mvɂn�m
ƞN��;�n�'�N�C�X�#Æ�U�چd��?]fP����c�\%Ev-,Em6�u(�*)����W7	n������N���'x���
jw�E���g��/�z�½�����!fE��U��b��r��+�+�e��N��GMQ(�[�GᲓ@o���aޱ��? #��=y�)�欿&����uK��Pe�=P�p?���Ajj`3�Cuw7�!�7�8��Jc̙Qe���|�t��z��V��Pa|�º�@1C+S�.n�%#$;P�`i�Y��.�k�?.��%+{��yMt ����;0}��)��yF��t�9z�	�Y���ʯ��3��Q�/4���YY%(?���X�+�V�W��	��	�7P�7F�Et�G��S�t��1Xr ].lb��v�����F��:P����.~�UDw��'h�@�<��ǧ�C�OR��LE;��K�u�|��)�@^c�\�rN�˩�4#X�����p����a��)o����p�u������@l��tN��;�w����
��r܃�ԣr.,ʻ�TXr҈�V����E�4D��h*�N�RF����#z��!T�k~)o��s��;�I��w�-*�R����������+v��X�Ry>0���+fq�����C6��g�*�(a�"^��BN�C��Li�4(��X���<HZ�U��#fA�e��IS�._w��5�|�	��p�j��^��7}S+�3�T�V�s����tI�'W|�����������#+����H��	�mGF�mq��b�@�ۀm9�ڳH��ؠ��!J}rS	�Е��[���a�5B-�6�o�y��{�o���������V��a��i�X��=�:' �b�	�WB�7�'�uN�f�Է�P�7���욏�S*��M�-�R�"�/�;��B��L��d9|�ř�=ӛ�6�CAĳX`p�k�
p�d;D��� v~�b�A��J�o#�'B��C�D��Y�f'����s&��;pI�� 
r�_��I�nD��shȡ�[eK���=�H�a�pU��ot�m�E.�g�(��$.CS�ߩ��N� *�����=Ͽ$��ۃ�F�m���f�� tO��R2�@���Oˌ�oNK�]�[1�:qz���+ϛ�N�2)��Hb�f4��jJ}��,�����<xf0���+CƟԄhi������Ww znf�������Ԍ�JR���*��*�W��%�2��pΎ��A�y_�G)���t�\:u-�evY?��l���xWF�ݚ8Tq;v���W3���$7f
g!�Ѩ�|FO%5%C�} ݆1U��4%��wt\����a�������Cy�����+�OU#���SM�;�:���v�uQ���)��,I0���ðxN2�sP�|�KOU��!����w��G$��@@���Q�.�}L.��f�%|��9v'E���s�&yf3.#L�?,��G�)��>���OӶϸ�d��a������!t�8�Z)������!�ɪt��;���z�5j3k��&[��M���m��^°u������#�E�����o�n��AJVy�
�$Ȳ1��o}dЛM�IP�~��c���ǘ�f��Z��;���m�|(���*�Zȫ�-�(6X��,g���H}�p�0L����Y�d1z>���z���!48��=��N�p�.Y��eֿ2�o���s:��ڰ(�Ule�x��;�� h�ި�6���zc�^�^���jx��" iIc�u���c"Y���e��E���?�h��S�V�<�˾3>�ڐ�I�Q�Y'͖��z?���:��ӷ��ht�7p������]q`19i�8�݃0@��	X��=(���c��0X��Nf2_���z?:'5�:�y�#eg5��O��'�f����5=H��sw��i����Z�����_��L���������L�0�� ����ቚ���!<3��b"z9��F\/^���7,�����$�(s��-��a���Q��2�I��(S�N�wX�W�D��v�RVw%�'!i5����U.m�dhgăn,x;qn�%��<Pό�Gq����q54�XY�����	v:t�cۧh.�1�0��5���f����{-b.o�Qy���*hu�ޮ�Q^��q���R:��8�[�̎��Ѥ1̑y���+x��s>�����"�1'��"�ۓ�G7���vv�!��a��"{��F�p_�	NWxy�E�M���A6L�zp��9I� �����}�����
e��)�f#L	t�o��4�t��eY�ڊ���,-�����v+\�Ch�E�/��§�����ߓ��ߥ��`�KRV-��ne�Ʊ̅#x��d	㨊Ih2����]?*ˀ}��]P��$*��a'��U
^H�׽t��B�gOR|#%-o���Ҿ�?��7ڨ.de�HK(�آ��d��q6�Aw�.�z�O7�s�IMf� (�&��i?��4��,:��hɿB[
0���l4�̠K�,6<��F;�y�x�HB����2g�$��h�,�8ZˋP�y
]�8�t�:̷�R'iO@��iB~���A��H���Ǡo��z�3��<�/��cO�{]L��P���y��Dj�8K���! �����k�E�y�9�nP��=rB1�	D�g\)��G��Y�^�O�v$��4��)�V�į����u���0><��D���H���@���Q������0F�����cIx��0(KT،�*�O�i��⼁�����\h�B�(j '��W�oA]+�Oo���Ũ����;#e2�ֿw]�/���R4]pwb�����!�/�H��? �{MG�xO���L�r�b<�L92�����#��O�1&.�5~�S�0�w��'en����X��xԗ�p���G��|��n#	,^���k��m�ث\f��ފ�J�s��+u��_W�w&��2a0)��=F#?���1��Q$/�J�$e��Op[/x���3����|=6�H�,����Y��#p�U�� "5�d�݅}��rv*��zx���*�#_m=��8^�^��R�0����EŒ�R��u�U��k�4������g����J��꒖�j�\���+�˕�+��_0��\�����=���%ۨwŃ~��t�@��jo/�,�8��[�������L)#ޙ���A�W�e�{��r���Gc�TP�~0ånz�T�[��A
�Z���|���v�]�Y���$�����7 ����.����
*��1P*.�.S���C�j��GUm����W3(�*O�Cz����2%�5�}��;���mdW]r���Փ
�>xS@��M��Oaz9����\J�̸�I�+(Z�v���D�t!<xÊ������ul�[R�݉rƘ{�K?�v2Օx(�:"|o{o�J;�HNN�+1qk�3�9�A�֔�1�������?�>����AB�Y�H����W��I>��s�J��į ��v�v���^J���:�e��M��/���w/�]:3�����+|6�������t;#諭�-��F��[nM�:�2���͛�?����X*\�Uf���xc(1�
��Q,�U�������	0A9)�TMa�N����y���T
��cY�/���}��V=\TDe���tV�����2���ʵ�mw{+��5�"'|*r�}Pa�%��L�sÛ��a�0����6+�Dt�H�@ؽ3��`<�@��x�n(!TP)�`�,Hgā �+����ۑ
6��U���K����i^�|��ЊÙ��&U�2��oU$��W�JC�`+�Ǵ#�$��@{C����>qI�G�d	�BRfi�)��i P,f]��L�']����a�M��.q.���"��L(s�I�.rfz�g�4�Į$L.SN�N�crd�&Ui����~�]�������EN{�|���9��u$f�sp��穧f8����c䈜��p$��w9fߢ7~_� �l9p�.���{�f6�,�.���wK�yYs����h�f��*<V'v2��iTW.��XRrü������2,�Tq�a�����Ei_�-v���b�.HΥ���7Q���k��^�	���KZ��.�b�	Rƛ�{q�z�HJ��g��B�o�u����0r�J%1V&�\漼s08k���K
c�$>����kRZ�%@?e�=��U�4M�rda�א����!��.����E�<�7�3��5�U)����1�`��.�~plp1y��G�i%6�������=����a��Х��B!���T��)�N��^�:�"����Q�J�M+[��]��E9��E��g�G>#��@ܩ�+�=�������`�BYm\4^P��@u�%�SW�Scw�g���S<���حU��;��m�a�l���F& ���B{�_G^�j�����k� �;�[�\�Gq�%3a	C�;����j4?7!NM�"|�����Mc�ښn�����#�(_r�_wo׿*��;2�y%g�%'�bэ�Ga��u��t�9�	`.�;��q:�e�� ��<T=��VG�>W~S�F��xlWM�Q�4M���u���	��p&��,�{v�/��?��	I�Y�<}�_���,�P�y\��E:�����j��w�ZNu�(�r�0n�J�c�G����O�R�����2��߅C~i�r�����1�w�tN1T�K3����X�D��)L�<��O7(�>�E!�8�5���v.�Ơ�!yC�|�i��M�s���kB#P�	�p���f��%����k*��l����Uk��!`����{��^e����a�CWQ��F�Q��lȣ�|�X��'�S}�Υ��In�!���g��3{��:n5h�%��("�����a��"����Xf�l!��jF]9��?+N]�;�l���w��6u�$
�Qj�u�y���j��כ�WN#���!�:(��ch r=�,�)��;�ڧf�rs���	�+��R�e|�aU�k�!��Ό��2�DK��> ~��l�V�A�Fc��qx�w8r�seD^�|%��N�.4 [��{���+�%��5�a,��g�\�NY^�U ��տ�C�dL;#-�����-M�ٰP��ΧH��QI;"�31+�XB%,#�Gaxڣ�;�h�RM���sV�QY�g�^~�f �=Gwg_��8|�*��lS����o�WE���W�?h� ��E˵����1� (T�)��΃��Fa	�k2ߎšq�����rO��tA���(Sks*�J4������˩����F�WF����В� �����x�"$"��Җ*�!@�>�����l��WP�B�W0�J�ޢR��mnt )�<;�[�n3�1���t�֬�5��B,����Ɇr�<��"���T�Y�
uގv`͐�裡�GƵ�"�>y:TX�mM����G�xBLWl
~��P�Лk+':�"�{�@��T��X"C�JW����^�r�ȯL��&GLnf�v:whA�{8{��|*$[��߳����ʓ`�{+\�>@���W�&���-%����{15]Q�<��@\�T�1Z����V~�7�B!��HQ��� (��oxv2ۼ�J8oY�Z6�=d��Ĝ-\c'�r|�K1t�|���Pjd㽲���\3߷Y%��jf�U��;�_@.�!<��Lh�L�F��1i�=����v�W,a>�fzc�Mg1:x��>��-���~�;��������r��9�] m�Xb�Q�.��+�
~����0�������yBH�uB�s���i�ޣg&1�"�@�dD@�1���p�3M`��P/�7���E7���T�����ˤ��9N��77A��+L�m%o������gG���G6���At&
 �S��0��w⩜�|/| �u�+��<3��RS�O��c�d\��,i/g�5*q٥�6n�OlQ_�V��<N��EtO��q���[W´�tܠ����n��5'�E�Z((+"� �ӾT)v���]Ⳬ	�I�M�8�ĺl��6
^��KT�~`tP���ELboȴ�w|�4�u0��kn�d��ߗi�YP��ϦC�h8v�_6�Uy�gM$]�	�A.!Bt�n�^�
N�f��K��t���r���Fߝrt�J2�g�{@�~"2���`Izp�o�c��՞SH��@~��5�|�,ٹ�Փ�=��?�S�^�`�@7lE�ƅ���#�p)#��*�����[��q������������ �O��7P8ДE�K�t{>��/NG���t���칏:U�h�\�M�
��2��8���osǐv�2�#�^@�r_�m�y���W&,DcQ�����}E�Td�w.=2
�y�U�^���wB:]�����h�&N�s��lV�P
�(��yJ5�����J98PQH��q�]�1AX7���3��Y�)�0g$z4m�l�DZ��G8����c�e��wO�m�)����v8
�e��6_h�� ��㶥���2K�!z,T9i�ךU�u@x��~�Kܱ	 p��=b�_}���m �G�Fm��p��+M�^�1ϔ���˕���	�S����@r+�]G�jSv�ϥ��Kp���P2R`�d�d�.K�TK<5)�.�Ȟ"�lq��hf:w�mKk����S�U�������M=����?Hq�Ӿ�{����K�*iRkE\#R�Z�D�
K�?	�:����/��%�i��Ѡ�ssx?�S��A��U �md�*�C"�h���X���%�s�f4�`�MXӪ_G^GR��2u��M٘�W�9Axc�&�X^;+0]�ғ���z�8\?�ID�7P���\�I���&C{�I�5pU��y湼�xS���O=L*D���c8ߏ��2��@dI�-_v4��	��!��o��zp��j#��}}1���Ac�a�OYI �$���U����[�9bXK!.	��b @&ge��H ���0���Wl:c�5jG��cr3��v��E�胆4Gc
#� 	�:PM픀ǝ���5��C����-�YE@�h�+K�
��i����%M9���m�#��בv|A��+�t� "�y�iD@-��!�+�Y����Z&EZ�F��N�w��,nkd*"^~Zb�L�;Y���4f#�f^�6��Q�&�b���k@gJlB��|{z���	t�����ˌ�0��S�i����W��.һ �Yq!�eO�`{��hn�>�N�G����CA�7�]�UH�&��w� Yʊb.N��w�z��T����'���ܬ;��W�����[�U�k�P��F�������.�[�����g%�8�H�FO��;>� -��
ƈ!m���'�x�����h��w0,�sF�$��䞇#���QH(� <X�ѿ&�(7n,�*Bi~�;�b�q� 9��$H�oh�g���Jɲ�wմk��<x6/Z'ɐ$ʌ;��'�u(9��U��<�~�������VdG�´�4���*����C����M���7y�S�֌�d�E�; >z�'YUF��А|�s�B�ݨ��̐�%�'z'�΂�T�^ښ�<��T��f?�+}���"�Bk�7�I���#'�������8���C�1[�z�]�S}Y��# $�Ԣ��k��h�����@W�; b�U��J�S���?0��J5Ou�$��b�u����/"!�?�_�� >�5����O]g7Tf�Yoꞑ���W����{���b�xJ��2�*_���ih�Z�
�$��w{�\�t]<X�o�VR��V�Os�x���8{aG��q������������A*�͌�(8��	��
@KR�p�[��\6�s�'�=�v��z*�"��B�� �X9
��_�?깛%�qO�Ԥ�;�>u��Q���V H�i�z��^�c �%S��5�~���/�K۲#�!�d�AI���>*��1��V��"�j�kF��U�_�36�m���-%�IA.�����'û�
/�f�2:ä���Ш7nK٪�]k������&$1�}����`�O����K�8�i���ߖD�"�vy!H?�		��S�y�EC�L��� �ېl��f��ۗ�-&��m�=��m�	�#�LLp����M�E0��3]Bp�d�݆�&D6:�<�>�h��И�o�A��ZH��Zr�?y�s���-�K�g�\?�.IlF�x7��<���o06u܊��IQjf�/.�f7�n {����pQ�K�7A�}&p�F^��|ֹZ}q�����
~�]���n�DC鈐���ꁚ�a�|�I�u�c��u����P3.� ��bv9� ��AL���7����Ov{^���r�O�u�'k�ް8PZ�t� j��(�LS��1x�!V�reg��%��9��e%���jh�ˏ�f���y7d��&b66�P5{�Ka�ӹ^+� g~��
ܶ����-Ԇ�U��.:m�q*�i�͠���5C�����^�*�Qga`%�0�&��Ka�V��5���]uV��͏V�W1]�ō��]T���@�-;{Q���lO�9l�r�6�vY`x�'��j�H2�7���D�uY��	k�Kj�03��Z������(�%=+r�b%!r��0��I�<g
���q�t�5x�IK/�`����~VB}��������N�V�wI`�l�-��8b�}��T*��e�6�k��u垓���Vi�e�Vѩ ���+g��sہn�7�v�/Zw#��ZB��+J_���`O�������+WN�_��8
{ót/������x!H�艪�3LC\տ�[�dp0��O��J��wP	2�ly�=벮��l=x��-Q��M^4���~!�[`��}�m�k����ץ條��lM�Hލ�Σa���Mm(5G"��#�@�퐗|��?�O-�	�	����|bM�o�V��H��p�(��^�m*�b�Q���8��_��Y���[m��O;5�:aW�����C�k+�ת��M��������z�����Y�2SJ	|K��CH/���{�,�E��� R��ûlP�3�$�.}$�몵2�����c�(��~�����aN��G�r�wחS��8KW��X��L��Z��*��F�/�_7%	wHI�d�γ"[�/ԧ�=k;����T�v+����@���hϑ���|�н�>=�ݕ2x0�2�1:�4- �S�=FO3]=��kk��B����|b��w.�pq�X\�q��/�3\�Т}(J�5.�)��G��鋲tJ���C^~w����{9��}�C�j��dS�2kv�e�K}��m6���|����/�J#��А�F���4,] ���s��*Ҟ���	���6����t�8�xgBUB)�ϺuRI^�Si\�FhgZ�3"7�J�g�� ��0��ձ�+�y����:�x�� "�2��ma�Zrr�@I�D_QF3Y$
J����R"~��E}lE�~���w����-��0�8ҿ����K�̿�K~���S�e,-bdL�44>�|g?�^S��30��J�&�8ރ��:o)}������ec>Kc@�.l)����|�mj)J|������76�53�J��0�r�u�r�82F��x����߬�@�9!5M$��9fƕt�>�������43H�(��4t/�Ck�D6�C0ODg�����M�ʡ͜�t�!(��zx��xB[E[m�������m�(�]��g��?��xZ1;v����q�z���ϼ�"�a�4e���8 G�I9�%��m��y �x&U{�w:��n��P%�u�!<W;��C+1j��?d� ����Y�:`$���!W'����Z�����,<m��4gt|,��f�\�j�n���k��,�;Z~��d�Y�O#���5VvE�ֱ*��1=�!�c,�D�F�s�Mܙ�c�1RB!Է��~v��V��b����C�#T�L�"=("���x���]�ՆH^ӑj��	����n���>��(�0d�DG�@C��a�ב�E?��}�6����M9X�H��I1�Xf�bٕ�x�Q�Cg&{�(,�]t��&�L%�Z��מ%�S�{�,>N�j/T*��e�mʑ��(,�^"��-��ǜ���������-�
�Y�X/{E�+�\-t�HGcq�'&+>27�;��8��O���n��+1�߬x{y���ډ��o1�4���GO]���h�*;�Cj�0u���u˨��c���*stVY��!�
�T�yz�Wx0sv��,����.��߁��G/�^�&�{C�w�������c/��Xl�����R�> u)s-��;��ا��^s^�8ԕ,�4͜����w �&�겮.:�?��qG2!/��)�t�=fo"n�d&&���A����Բ$'��;&?�v�Q�j�ǖe7f���/,������@XǗ ��o& \ ��& ��?�C$8Y8���9͔�|�K�VȾ1�@�x:�H�>�4�Z5�W��ͷn�&i�Z����â��Z�%���E�*Uh��k"���su W��f�g ����+�Ж�So��W�=kSb R�7�2���:;T[��Op��Տ��P	�p2$w�*O��/�#��@��[o1�)#Y`�[��3��������/�������r{2������(P�9"
h|���g��h����8�y�Z�Ѹr��@���E`U4�S�<�;�u(�݃k����&�6�ͭ����H�Pv.
�|c���׌��;�(�)f"jq��{�~L�J��<���HS �<�"OmY��ﰪ<���0�!6�{����H����Q �Cn�"E���~���5p���Q��vF�� �1�q�)Y(��M�UQJa�_����S�Cu��7뭬���SY��
�.2E�8Ugc��eMɦ��'�cJD��[��[���ϋ��`u��
������ �\U#�6U�c��?5I[Ȁ�X�9B�����v����aEInp����<_X��dĽ&Y�_jI6�GZN���\����aJK�3Cl^䔯�+n !7V�ٱ{V�
�� ����U�gHv�
��+��٠���Z�Mc��P�_��.������R��&�.�ͳ}LE���
�}����tG�\Z��A��6��J@;y�J~p�e�BVb�0�cD���F�9U�F��s9�5�6T��ñW�=����~����� :���!���n�i�J�*�S�ͳ�(�Sp�&�Ή�-\W+߹���r�.���CE��,�48���î���c�]Nu��;+��@v�kW��O�e�}ܹ�+=�1���δ��U��Y�ۋ��KwJ�-E]�0�yw��0O&$r���^պ�En�U�aD3.��&����X�Q#P)����^��r�춦�e�Rcfr(�����V�ֹ�� A�����D�S�im���dh2��C �E��9/�ѥ�cz$���dg���S]U)���Q�&�{��[�3�f�7p�Zw�/�� ;!g鱩֫\v��iB�(��%����Ώ�
	�x2��\��"�6��f05Ɛu��U���w���$�\����{�9,�؎�/{�x��e�x�����Ъ����@����*�Fi��3s��J�K����-��]���YZ$-�5�4�G�D��
s�j&�cC�"1���)�Xم���_���'��y-�du��/���.��*Kտx�}{�D�n3U���+�;��ީ��z���'��<M���o�/)!���bھ�q��dm���?R��W�a�#�6a*�x�D8^�񔤎�b~�j[J�v>_�E�Lw@4�-́	o���e=Se@���]���`�.+�đh�ϫ>)�@�h_���n[H5�aԲY5�5�HV��Rǫ^���	�Q̋��m!�1Q�q�;�+��cE�C/P�bT?+&n?6T��wސn	#$�"�1�̬�Z����o%
8̬�X�;��� � ;Y��gl�[x�m?��\��n�K0�TK7����،Xp��g��]���[B��X�E��5��7����MZL\B�Ⱦ=�V����Mny�D#�});c˵�C"~�C�E6:ɨd,�| ��y��8�	�uh�p�H��6�t�cOjwm={�L�^��*�} HM�q�uj�C�J�	L��LN 1��p�̿O��{�s�~ϣ�c^�}��H��뢧�^RMg����VrEW�p�E=�����p% ��jr�*���w�:�v�.��7ٻ���C�u�rb��ӱ�*֖s^���`����(�_!�/2h/�s��7�����|���,�<1�d�B���`�%͜k[U��*j|8a�ͺ·X�V���dh� ��F�pl%$)����	)+a����c�;X�6�G����{:�m�]�!2/���O�ثa���ܠ��]�wb�N�Dt�Pʓ ����&�M~�I��S�p�P}s�[&Ͷ��^G����(]���Jã�י��U	zꩡ��u�ꜝ� ۩�뀽G�O�.���*:�=|.�?�Fg�L��т�˭?Eoi���M��~�6��)���V\�	c�D��Q��<�%&��3i_�)�I�TQ�D'����+���
�<,�����ܪ�s\t=�\��ȦKrˡQð�%9d�B�L��jġ��/+��;ƧހZ��K?�Ew� ���f�N���,pj�YY��ЦW��笧��Hv#�;�Z�&ג�*�G��{Y�x;�.�§2�������<��%��7���[ �s��7h�t�KQ5�k� A��T�?� J'T(�c��������i�i~�l���@����՗6����|�$�l����|_{��z_�3m�������8�Qp�h�
����#,x��+츍~�5�ʺ2w�κ�/�I�t��G]�pvb��{�g;J�2�Wl��B{��H��v�v�[�)^)�����M��Oy�<8k\����x�*���&m؂c��LW��k�	R�.�W��v]U�¼�e��ȋ]�OkE��?,>V�J[҆��q�"��K��׌�OC��RX8O]]��a��H����6�J�uqFr���Y��E��"K>��+#�U��_��H�qYR�F~[��n��d���lmU�i�=v�G�l�U瘜��`�V�Oz����a�e��e�Dz�^���,��B��
}ț�0db@+�`ƀ��Q�RgS��.)�\�·���'�f��(�0�XLN����1orPf����!*9��YDz��s��y��F���صI^k;��r������F[� >���ty�v�a��-�A�b�݉�tV�,����E0=�/ﯠ���U��EY"!y����L*�Lo
Z�������P2ϟO^gW��z��w�n�����R`n0MyLkU�0]	?b	q����{��Y�euU[��2�b�/S�68f�x��V ib��yc8�uo�|�UF�-�ZU
Nn�М�4?ھ�D	�n���fZ��歎����e��(5=��ɚԡej���H��&A���ZVL�0��^2G��V/�{ǞN���0�.��OT�U�튥'���g�-/�r���fDq�u5thXp?W3î]~Y{9��{�堈O��ϗi<�kweLnmx��T�yG*�������mt�\
�>�)�/^�}�w���W8'���,�)�;D�R�($�l�u���D��VL�-���}����<u�2�e���Ys���[���kv0n@x���Z`y�_�����G�=���j���_/��^:.`!`V�s�X���i�D�ó)Y&���W���-L�T��Cn�S�K��|�-�J�Sx����M������?����T�ϯ��\�{J��I(`�j��<���(P(��)��t�4ĝ��]�q}e1�j�2��؜�7�a�d��I�F,�2����'����D�R,+��i����)��#f!,�P�qQ/5fp{ld@�f����"�Ηr�K���J���8�bd!OޜT�q�Tz��B���e��k�wA}��+׊�S(�nA�Oj�
�0'��\�j@>>��f�̊��.U���`M%�\�̕ړ-b�i�[*=��ӡMS��c�8�.�����,Q��5?�i^y��:y�n(54n�H��m�o��s�(HDnXۍg�T�&��8?�9��Ҧ_�v�a�A_!�Bi<���-j������
l���_��?�)��v���D�2_H�:� _U�Z��ϋ&���N"�wO�}�������h��{5�E{�\W�W�;)���y�@䣺&"�%������`�Pi��$�o̠��������`xp/~��	衋x����J�.Ǳ��@1����x���6<+Qn�W6�x�ʹ�~�S���L��L�{ ��+��s�H�U0TE~$|0-=�j�r��IQ�lA���>=��Oo�С���P�^��,�x^�o9�� �����i���A,��������������Ԁ=�,a|��}tN�!m��]W)������٬k'O]��p�L��`r~�1�0_@�6, ��1n��T:��B�۸ʛ\͙�ڥ:A3ϸ���8��O�SW��1�䖒6.E��as+�]�vz��B�K{!x9v����� <;���qn@�4谈��@ťP�Y��M|�/.�K[��4�M�y|���].��E�JW���8�4a�t� v�d�C�D[كQ��,XJ�аu�	���[Z�T�����?�a�=���!��G��C]pObr��:�?O�ymP��ʜ|b�5���^�b� �uw�b�#�r�Y�ߗ(&m6*�%���X�8�"�xB���O<�0F��nL����m�4��\!�������|�6.���k�����Ϸ!�U�+�� ���R�W=�I�[,{ڮ�;t]P��O�Ċ�)���6 z|��m.8n�vCB׃(�;d	!�:!������3�i�"Kά�&-k����d��:v��+)m{�k	!<���R�����E(B`�ۚ�hWrm���,4��_��j��韴c��� r�a_B���f�O~�����N�rx�ARUؾ�����`?I �쏤+�/�lIFǌ�N�)�I8�:U0�.�BE.� ?�&Ċ��o;q[Bw뤂����-�j��m 9��^ɿ�ǘma�W��(�A����16{c�7���g9L5��nqe��%�}J����?��:F���4�m�~�9S�91�Θ7�Ӧ�t����N$>r�W:�Rj��'�����pi�^�����R��l~�:˄�>H��h?���������`���'��M&���lS9�Ѐh5Њc+t���*�IC��.��k��"��6y~�;?�]G���"����_�ja���ql�e��0���.!��Z���.�l|����sz_�0����C��h���$��cQ.!	C�V�7s�	�#?K��k@��{��B�_~��R�$����ͧ$�u��뤦��&�}�n�!���l%J�$��9#끮$8e��^͚N�%�>��T�x�Sv\����"[�#����r�xvc��^���:z���q}����EO��'� �Q=���DAݮ
7���{����ލ�+�xE�����X.�Wdh�����QY>P�����ݚ�}L�H��h����q�TMz$qm���O���n�����Ȫ7���BET�ꘖc]�&��;�D}6�!����[Xw�/j�]M��7�=.Q9�}x37�)�� <B)7�չ3�և }YYW��=�(&��]�z��g~�"h�I4@�#I���|�fۍ���p0@;&�s�Inoߊ=�9Q\V�t�b��Hg?P��\�:�Gؖ�o8y�	O��;2<������v��]����ݎ�}�,����$�AE�����F�Ǎ6�	�8���Y�:�������J�xH�[&��ejkzvf�\���g�7~��3�D-B8;��j	�ZN��
�,=�t*�Oy�g�r���NI�(g��I�J����-V��F�7��dK�2�����,Zş4����5#�_��6F�Dw�[��ո`��E� l{�R�8�̣d_���4��r�����wN
Od����n��[g�[5N9��vyb���u�`Ǉݩ~ )���bS�ˀ�w����^�������8u���J�A��b��y0~�qIP-�fN�TJV�BA3KM�6�JeVU|x����ج��2ʓ�v����e�`)�F�ہǐ����:����=ф��:��`�v/�0�?�,!ŗ��s�E��7�kȕn{τ~H1�%�b�bCvˡ�#��v8����������4)'G�=Y����(�Ւ3�A��>|[(15ɼ�ݮ&�*�1�.'s��XO����!葉�ph�r# )�������j�@�r��ˊ�&��H���3D���I�}�U4o�������!���[��}3�,�;i�K�.����G�F�>Wꒆ�Fß��$/A _	?���3fiU~��S���E]����M�O�Cs;b��h�W�/Rzu�����H3���������^Zu7��z^��s����5L`q�U!ՂtF��o�pyj��b�Eح�ǳ��x�I��<��,�#Ŵ��(�]�������I�2�f�tɫ�}���̽�"T��$E�3��Ѕ��S�|�*�d��뼊�k0	�f�kvߋ�>l?��X�`S�{�,,�� �~��iဒ��X�����r }t�H�ؖ��������:s���@��Qkt��\�2���`�n{i�!M��C�+Z�-�8��C�vKޮ,)�2�w���Eܠ���y��|�u�(FQ2�F�E�@6>��Q#��l��ހ���6�m���c���C;w�n�7�*�}�J���n�Y�Od{�x(i�\ht��� ���Ǩ�\"���]���Wው�pF��4X-u�2PL�~����M"��)��m�a���٦{��� �yˣnK` �:w���jX9��;�]�5%���~�|v��q*Rm'�f��K,{��b(d` 9��E�؏��J�m�*W[q1�b>F��}����]����&lQyY4����-Rz �!L1�0fA���u�?��1e���v3�E���9+��?G=�1��^�A+�b.��$���rFqv��ª��a��WJbL�҉�c�k�P�P��:���^���_��V0��`�B�Ta�j?���$F����[o/^���a.��;8m��eG7,�����D����,Q�b4�X�]���`|��tN#��g����hq�k�������]��A)N �93s� ��_�J��(�B&{r�I����	���tb���	{P_�C%����2��}�!�m�H��c}Md�^'�������>�|NJ����Ta�ʉ2��J�q��޳jz��������Z��u}�����H�:�ҩ�I"�.ݭZv�Q�l�]L᪠l1��>���͉Ԉ����t�ǀ)�7W�sY�S�ZaD'��£xX�M<ɡ]��~f��ǭ���2�V:oV�l��4���Kr�F�Xf$��.P\y�����#f���A��
�VP�&t��-���5���ډ����R$Z��N����,��8[�{��`�!hͅ�N�P֦�8��/d�nX��4���#n��@	S�S$�mڀ!�c��_��o��\H")�,S;����p0��oʸ� 4M��,
����4^hDp�A<��`�y�
��,c0l��M*��;*�쁄�\(T��}kl���r���+ �q���o~�^�Q3�jBxBp� ւ�ϒ�.@ǐ�ǫ眖=n�mcgR�t�^������� e�ƃ���*N.�����%����y��C������T������^���#�hm�fS�XZĀ�ݘӓ�_��X�L�����!�����Q�CAK��k��J�uNѕ󐵴Q$x�D���$���R^��!ԋ`�X�#!�aCTJ�VE���4�J�s���w���E��Pkha�%�Dn�_��0����4��#T��UP.�$NlD�w}�)�zsޭ�ʤ�d�3���
�2 �E��@ؐ#n���Z���3�4(pYvVA�&�(?D2ե�����%w������$#��lɡ�:83�O��2� �����p���ݗr����{e@����E���	�N���V!��6"�6��eY� Da�X����mo�B���!�=^)��ɠ��g���\r�Q�gp.Jm�}��e���e�Bw���۽�7^��T/]z\�����438$F���t��1��/�I��$������ao}	��^�um��4`�"�-�~}�׶u��n�+��X�_�U�ĥ�AA�:4��DO�b!�B�L;�;%���-[+Y�ɋ���
���S�9iJ/<�:q�C��28MΫ�Z�y�1Z���'�����[N�� R���2��|�o:(�
3�	�=�n�jK��O9�t����ff�����y�@�Pm����~�(�
�b#�.�y��'��<j���7J��������٬��9'���q�fn+���7N^�D�;��m���e�Q56:>V'1�T+-��V���;V��ŊQ���uL���|x���x�Mi���Q2�7��%�/!��],�YV��>5�I�t���0��t�J�j�DV�8  �a�-_S�$�.��D��@n`����uq)!�/Vx7H�հ�A��"m;PCd� ĭ؜l��X���ع��/CYH�h�������kG&:!Lέ�z���M�/
���R~�E6�J��r����ܿU6�ī���\s���R�Ir��T����#���x۶��!I�?��=�#~,u����[�c�z�1P����3��8v۵n��39�`�(+Up[���͕EQD6������"��#q�Ӕ����v�$c���Y���yVJ�1~�@���A+ep��V3��LHϝ��9��l<�܄��姽=��"@�?a�����O��z�T���=��@��(XΫh�J��[�<;��n�%ЗR5Q���d*�S�����0ؒP9�,��hL���A1�5GZ�?V�2NxdD��t&k�Q
�Ü�qR��͛��Ij-.����5I���*������ ��-x#��I���f:���'n����8�����2�x�;���Z(犂X :����ϰƖ]���Eotx��Ω��q���lbT ,�h=�5M���P|���g!�r6,�,�j��ﯳ�=�g<�����~S�"q�u���"����k��"�6�tX�y��h?�D���� �����n�M����~��k㧫��^[v�r�Q])�3x����G�-�����ɶ�,��E�]��)(8	�`ő^x[+D|C"�QA����h�NC�f�:��0��I����KX���Ӂ�%�������դ�����D�VK{38�v�ŵo��$�����u��.5���g�\=�T&dw0������/;�됩!�
���>��p#�@�3��_�N�`�P�������o�y�D1t��G�����3I�t�6���<��Q��7B�{��qm�3�_4i��3����}'%Z����KOͺb�{�������?������~�����h ��d|e,������5�q]�i("�hOTW_���i�Y�|?�Q�3�V��7'�Io�n�!@���/ȣ8Z�9g*x:����6:��:���<4������c�x� �8����l��ʋyM[XZ!-++PD��$Fk!�A&�j���e��&*��;_��+�'X�����h�2��\��=
�}�eu':�Ì�tK�������(�_n���)ڼ� �Ya��T���+�[��7��)t��"A�UX�4{E��-����Zk�p>��e�v�E�#��8� ]���H�-՜O����6��b�+OKp2x��<k(h,�;�ޅV]�}���˓���e�)�E�{h�>a�e0���[�M�<����~�;�|J0j�6XW��2+6�[ý����$��J� ����X���\�7L-�n_�./��� �p��V��ZMs��fz\v������#���6m��ɹ��i=!X���υYA�o��z��i�O^?�$<Ha�,�d�u����sm�E�	R����^3{�It�@k{m���� �@0�~��9��E��	�`���=��Qug�u!�f%��62@���3�:���={��GW� }4 �+)y2�p�
칶��<��~�4,��Q{X�-��7���\4�z�x�)P���l�����lfAl�����c���Լ�_%	���f��22(G��H�qjG2S�㋗ָ�	[���&Lv�ϼ>y���C<�ʦ�K��;�e�t�r��{ŵ��!�}�Ss�1��R��N��Ԧ��H����.�`��E��fÍ(�0ߩ����l)\�_������8��`R� ��*�	gˆ����5�*�/Zt<��jʊ!v�d׿�l�|�O���}IXE��0"���ԝ��k {N�v�}�t�����1��O���O����o����Ņ���a��н�k��|`�p0|z�iJ�	�[I'l��l�J	� �H��'�4�?��5y��S)bצ�$t�Q z��$.������ρ����H�k5l�J�����]
�<�u�@}�(�������?�5{I�*t��"�8�����G>��O�2��\:u�Ut]�H��7E�����z����p8n[����ŀ�Wn=����N���8�,yƁ%u���
l�E��M�����+���p��En�+1�nI�e���f�W�gyG��E2(�/�3�Til�&����:u�5Q@%����k��_�8:ۂ�NN��<�H7��"��$�*T������Y^7�\��O�e��vLC�Q�5́����9��Ay	�)�'�g��KY!;T~�]�U��~F� |2.lCon�J�u��֍jU@�����i��[]*U�4�J��f�q:/��9yha�Lzh�T9��#9K����ЯI(`��$��$�f����^�S�v����y��4+�1=ӗ�2�V�F ����r
�������x����AH�oDb�|f;��4�+�:�y�[����o�r^+{��x�4�l���@|�����*��.�C8jY��S��i��(�T�nG��/���ZT	ZT��*��+CF�b�r�l]LHp��>ED)�75�(I�Sk0X�3��$clי,BU[��YEE�ҟ�T*_E�� G7�W|��N��: ��T_P09���f1��C��$�"?w����$P�򁔏#d�mG�쏱�� W{�����	3ӣ�#�Ӈ[{"����E��9p]�e��a�D����_r�
��W�c%��� e��\$e�4��&p0c��*��S����q�Q~��ɸMw��3�p_T�i|�+��*5ά���}�*҅p�(4{���(�����/��'"X܌C�u�҉���1�V!�� E�j��� �����5P[NW�L��.eA���o]�Bd&]�n�>�A�d�k�z��u϶�&H�}�Q>��0��(|T�U"�Pt��P~���hU���U�����;6��~�{ �?�F�W.tE�>s�V�J���[��B ?�k�9�܃�+ff!Ȭ5iS[|�����W�HZ� ����;�8��'�Ƣ��4�Zo���Ö���d��� ���H'������RC�S��?���+Ǉ�us�]Y���-�A'2№.ꃚ�&���	�w]��7@���3�9�9O���RO �/ �B^��Os� "�r��Lx|M���'�Y1YM�4�o�������l����G������F��;�2�D+!���5�S��.�yv]�q'NPu~�R�d��Jה� Bu��،)������C��6L�B� ��D��u{��B{���}�x�M��/>ר�>;'��=>���8'���A�=$ͪ!���v�*V�r��t<��Rk>�]H�Wc���τ��"R�g�%�
bU�mMs���UU7��	�Da�/���n�L*���"8��.�-G� y�����>��~�c���b$��UL�E�ͻ�e8�1WZm쐄�}��ee(E��g\i���OZ'�\��g叇��5�2C�''����%�(�@F���ֺ��*��c�&G���� <�;u�� A�+�r�G��E�]m�y���2�`���B]}Yb�<�������XQ%��x�T��k��f\�����5������n�,�S<(��7��8��Y�eS��Ɇ�Hf���@H��p?���n ����-��O>]�d�ڶ��c!���F� ���Dl��-ͽ�!������Tr�ؼ��95��oIn������Cn�n4��P�?����Z����\�C=v�=�V�<���
ƛ�i�#����U~d@S[|m�����;��������a`��hǖihH�)G۝>�K��d+�����	��$#��ٮp}�e�؆_D+@*y�2��k�x*f�7���)�KE4}P<��`��3�Lğ7�h��8I��I�c!g�I�`����]��
���5_r�V�F�c�~J�!�@�=�b�y��I���͆�4B��0�I�z���X�J����W�{,p�^�ͫum�лiP�X�Q�A���Đ�y�译ܳn<��8�9=��{�^��Ha L >9����#�Y�?F���^�gr��<���('�i��}ͷ��7�28�E���2Uu�S�;�r�� �׶�+���u�u��5.o� ��(���5܉bD}7��ګ�(�㈞e����G��$?�4e��3�[řc��3��9�C�x��Q;�c��&g0o�]�4�Zy�vm5yh�j��c�u���o`�;�l�s��01ɠ�"����,�Ϋh=$*��{����,��,q���.��	���3T%^�_�������� jX1b �)��}�(j1�7��k�h5C���S���`�'�Q;�s hߙ�{cr�}d�i�k����]��]�M	��yb���;�yq{,怷�8��?ߍ�JH)�m	�ky�����x__������/W����������ۙ�b�kNf����e�,� %j�|��<�N��b��y���-��9$�~�r�޴M^�x4�n�^���'e��7jnvLC�����n�U��(@^Q<r��q(�CD&��W�cK���g��V~%�u
sQ<�.�x�h�����JA��ن̂�ɿ'������.�(Xc�0�K��\9�PF] 4�3���)�<t,yUG ��6jH�p��8�(s.�o�y�Ԟz!�W�q�y)�+�{n�-(�e(��v�50��H��fƿ]<r���a��B���?��r��{#� �b���ݠط�
T�Bʞ����S��0ZP��{� �_:2�A���m�~��#�������h;r�F�i8�����z�+ފ��I�I�{��S8��_�n�L��fT��:��s��q��|O���LYO��{�O>�˄�C{�=���ȅ�F�IGfX�#�}46~t%�%��[�F{:���"�9W�$,B(L�><�y�5�@Ý������@l��BE4�>��PnG9��PpU�:�ו�}Ê89!Ҟ<�odm^���2���m�>�i�vOϱMd�(�C����?�o�b��C�!Ր�
Y����h�0 V����+Xf~�����R:�41�2�0Y���#�b�x�Axe,��ٿ���F<�f �$r����U�"��$R2��~�Tv\ !�(�$�Zm�	�@	��Q��V�|s8D�9��  HԊUe���s[�'��{���-�W�|{t|��3ne�7�5ML��RSO,ȒWo�e�:Ç�:�r3*��#-�5��Q�<�ڤb�{�N�3h	��y.�s}�fN���TN/5}��&� %��]���T�B6e�s� �}�F	�ĝ�;�����[U�{9.�}�!8�w@!����t��I��[�]�WԒ� �}ר��,�b^
:�Z��n+#�<;R%�G⣕��U��K��oH���%>7���~2�ߐ�4�Jz�;U��k��g�ouQ?��J�m�!X�Hi��F��a�O����p�>�h���!̗,��LB�c���r��t�{����s���Y~g,�w���Q���!L3��c+�Wc�5�eϫ@ݼ�uۂ�EB�ʺլ޵UNQ��`ʄ� �π�� �Q FU\�|w�zn�
y���ȩ��xc� �l���k��b��>��@��6f�snU[�D�i���u��'F�n[���k~&[�^\f�菲º��N�O.#�"�����h�fn3$��z_Z�"�[=�mԇ0�XU�e��b�&d����'=���.8��'��*$N��\%C�Lq��p��%�T�*��^�t7�t��$�e,�[N���"6��I�j.beH�V&%W�C�3Sf���q���L�4�Z.ȥ�+)�B�4l ��@���A�q����)���<���XW�rX�*��(�u�������1��Q���v
;�/�>��<���Y`�p2|� �M�
x�8Ga+�� >�yg�O�c$�:�����v3�)�
�����mK�T>2�P�ȈF�]��vW�V&�o>D���_��^mр�(G�nJ7QP<�F��=)�I`f��IĔ���ߍDn�S�'�O
� �Ŧ���K�L�J�i#���P��c؋ ]B$eM��cH��f$����VJ�:�-"�0�7xf�����Ky6�TI���DĺR�D5�8��;>�Vr%�H���?�?��A ��gʵ�[&����=���ո\����:*�6b�*�-����m���@��*V�+�Y�f�u����GC�%�x
��&y�WeH�v�CG�;r�������`�k��ks�k��#�ތ݉��p���~�@p��z=}~�!=����F�lU�v.�do~���W����˦��	5����\E���)=v熯���� ^Q憓��[Ӕ_�P7Ӥ��E�D����E���得;�405Xk�`'a���H�����f���db�,f�AN`��P�HN�����L#" $�K��9Hx�+�����[_��7x�F5����`�P�rA� .ٱL�J��~N�j��b�,���7��ո."��+7ݘ�o__���Ѽ�堞O���%�oS��7ȑ��ǳq��h��'�*�m1W�P���U�q�@僚��V�_��%���mx�a�?C�Pﱬ6�ܝS�"����1|��{�Uwuz���@N�qd�E\�K	��L
E�J��}����h���l�+�	��&�P��ZR��=�o�����~��]q�SP�GM�5X��+b��螯*�`2�w����O�����M��{��-5�6��Y������Ќ�� Q�|גp�|ou��ڶU7�y��X�i0rt��pg9Խg�k�iH�{#P(�}�����6�������E���}+�Z9'v���S�yO¦�����x6��\C�H�<�f��9I�0 �����u$-+���4a�A( � �hof�.Zn��܂o�c鳺t
+��+��Fo����ئ�C*��Q���w��)h�+��v�~6�p����X3���Ԝ19���;�5� �Ռ�)��w��4��W⧶��׼�`}����08�p�B��~=�=�x�^��ѣaFag�L0�0~xO58m�x�_KbN���&�K#w�#�-N���N��	�\M���EȮ�X�)�=`�e������g�����\v�h�q+�|q�Ҍ�{|����xs���(�PZ�t_�}G�����R�{'"^�e�|.���]��x&i���ۗ����I���b��^�@䵬��(�(W�Ѧ��[@��<).�נ:O������5�M�����0��J����v�^���B�JI?3ƾT����1�)����\@fk�y�ȗ�&�U�>6�L�4��� ,w��
D�S��˟N�5xg�j�#
u��k�f�N�T�͂[��������HH݉��/j�po%�(&�fqq��*p�}ւ7c͏�S�2E�V��CJ�G!��0����L���v�r>|�����0���q��=���	ʙ�����.@���z~����'{mN�y���$�Җu������^ɼT!`��.�P��=5:	����utM�k�����CM�3���n�:�G�(�[ ��Z�h��e�_��xل���Ҭzjx�:�˺c�.���[�������I/u�E�G�A��C����Y�^R���]o�j��B;<Q�� ����c$�5�Ǽ��e�37��N��]C=�ٱ4Kre��LG~�&�y��Ȅ�2����C���ܖk�!"�a<��?sխ��%Z�фҚD�����IYa=.hmˀM��iP�p�>T�f����-�/o�\�?�4�8�-`34�NRJ��)q��Q���r,f��b��T��FxL5����YA�u����g��.�CXZ�#��Ůg��)R:?i�/�q��)?�.�c�AYR���	Qw̓�V�\4vX�.89e��)�E�c�ʶ[�-l["<��qr��Tx����GRT�f�xԁ�DK
�}��`��[5���z)o��"R��_*�F_c��i7�ic�Cs�fVHx��z(ӳ'IT4&�5��+�V���G���C�x�	ޔ�:��p�G�{�:e$��@V�3,������"��U�-n�������Gd����7�����p�6ei8���;x-�[��dj�?�~�q�F_��|� ܼ��y���\v�'�ex�!i*|=<�n%�kvAS�g��-"�Kh)T%s�>9zñ���R�=�VIE�>���:x�Z-��=v�)��U��t���x��h���j�Z�_BLU����B.���ȏ��0��T3~��\`͙x�12�vB�Bp�_#����#4 �4�b������}��(H9dYՅ[��uJz">#���;4�=x��?�S˯�������!=c� ����J�Dr^��br�x�����u�{$��B��Nq��:�SHS{~�<G��3I�YQn�h�����Q�N8/y'bri$�B/���7�2?���N�
��"ӻ"�	��gr>3���U՞�~��L�_��CTS�"K"�]M�O7L�鹝�P�?X�~1
��Æ2b��"?<�2n6�3��(�ٵ���z1�غ+��(u�#��p,P�{8���o�w�T80�`��G=�֛��XE�s1�b�;H�I�#�<a��{=?G-�k3�V+�q^��P��#o���J����~�+�_#Q�K���6 ���6%�pH1�^��b�� �m2������8���,G�b�２�wi��NX����]K+9v�����l�?T<�+��c`����-�+�`���d��=���ri:����(^���_���=%dߐ�@�EjmHN�cgV����{#+�,��7\wƜ�.S.8���B�	O������1�t3{V2픀�wbX�N�i�C*�LL�!�N�X��P\Նvs��n�r[�F.g#C[Q�ڃ��o��1 i@OK*�k�8y�����{A�sV�b�0�z.���oP2=�EGp!�w��4�Rx��2z:��P%���E.�c��2�:�3�]C<,��vj �ID��t���- �M�Q�������~o���BB�� �փ�0�1�"�8�ŏ�m��y��2Jړ�%<*-��jQ��0�f�
u1̤�;�o��ѮG����J�G�VbS�\6��<�Z�@d�RP?km=�x!��6�v\]"F��l��	'��:��6��K. 2��c"�}�+�N~S�����5c����t��$�4���'�h�5�h�h`]ue�ľ�Z\Y�����+�ฑo&�T���Q���<b	���柭�\S�L���:��n��GJ<\TKk֥J�;�Oō9Q;Z�\^���`u�@�y��;�L��.����������c%��-�U�!	�$M������ صXמ�q[�n`H,T��T.�9Zs��-���9@�뭘�@\�|_�∶l�H��,���f	V|��^k�ꔴ|�TH�jY���l}�F3��f�|2���,3vP�f\n�X���(�BV�8F���66���2]5I��fe	�-�V����z&�3A�)��8F)��Śx�^��	&�֮��|������ہ���7�����?D�J3��f�Ru�4�B6�q6�1+r���&$�|��>�o�(������َ�ZS��p�ɉѲIF���J%�ѭb�2_`ټf��#H�-v���ne�Lz4��wO����ś��Z{h�p����hUb�q���Īժ/�c,�C��b?����p�kLV����z|�j?T^�BJS��APv��sYn�j��,�*d%|�x�f���H�0��v��=+��BzݛP���L�Ɔz ]�E��-�r�͹����� ʁ�t\�9?#?���+C��0�}��u���/Z�m���^Y���c�f3�zkZSL��`(�;8�j��c\�{�5�j����Z��v�� f�.d}�;D�{�a��|��&s9�Xnu�h"*`ٵ�+�vA�{�?ă�L�V"�,��T�oTT�$���0�����^:'������혊�)��m����⃶>�����UV�1�CAm���,g�,�,L6k�3\���!�QST��$�c̛�n@��jxbP��7��12���.l�A��Ш�[.�����Ҷ��T�?���ff@�A��ʌ�2ن�i��c>3�F�U�p�W����f�4�Y-�)��'�b����U�<���.���'q�t��!\�8\�tS�F�m���'`Z��t����n�ҁC}������g#�_N���$@
�>M�3����r���7K�y�V?�������$`5Gㅒ��J�x�z�[��G!h��T�Z�ͽ<4��F��oj���?��J���	)�2pCa�%'J{����)�O
N��ܩ��|����P{�*���U؁�A���.0O����Wu[."���PJ�M~����'݃�ˬ��Y�B�
y��E�����z�D5L�bYW�(�i��Ǐ��<igq��W��:���B�Ә��K�*� ��?�"�4�Eзj����=\�T�K^��KL���,j�u�>��0�_Ch`��ݪ��K�_cۘэ�x�+Dx{RzF�����rL���˸�Jܝ�!fEW����[+o��Xp��:���5�O��e�[�7��ƨ��X�Y=5E���*
�s��03�w)�P�u-P����dt1PI:ֽ;1��L;�2h�Z1ǉ�YL����sSL��5��ͽR���N�ܥ����F��^bť�f Y4�?��8��d�+��c+��7���R��;*(yz�]v�[ͅ�lw�CQr���j#M!sl9���@M�9�_AE��VfC������%���:dzs��D�Sڈ'����_	E�ܬI��k���jC�k~4�#HQ�	�X_��� ��S�F���\p%�nEoՎ+��J\llIǉ\p�&����q(�w}¾��T��H̫3|#/��	�1��}� S��fes����k��5>���ջ�ձec���[�\a6vn��~�ʔ=�_�[j������ ���	�1*MM�^����W�8�"j�57rr������l��)��z���5f.�s�����5��Иz�K�<	�V��η��3fE�bl����A[����lۓAHU(g3�kF� &9���P��A�W���L�d�OeW
�\n�������,{�"d�n���.�����2�h��+�*6�-��"~�k�8�5R�6T�I�=̢��n$I:�؟#��=�Y�ʈLBͧ�&�?�,���L���Ȱ@�b@�K��lտ�*��ѣws�����^�v2�Si��~A���rdo�ĩѱ��Rw���O~x?[�����I��NI��yU!
��!2����#A:�_1��ZN2]�:�VG��Y�v	���z}
���⧃�
:���$��I��.knL�x/}�Bvw�=g.�����X!z�̡�2�k�G[	����qh����3��J
l���J����hm43�E-�Puݯ�A��H���Dk��Hl�ǈ)@n�ݨ�5���K��{=��v����ԍR)�W0K@�	0o�}/��΍��G�A(�ˬ2��/_�����L����%�ϛ�w���Wr�	�g�! ������L���&c4�x��B�}*��i�T_�h_ʯI�ٻȋ���F@c9jcq����]4S	�|�.��0�jR��A,?� �rt=ڔ�~�Ѓ� ���>Τ�[�ET��4ف�������Vfӑ���C��"�5�{[�:��$����evC�@�b��F��EåBuI4�Oqq��p+�˻�
�8o�;����s�x�X�c����7;����B� ���}N~R�y����L��4�֤D5���ֳ�4:�Ì��Pv�L��V|eT�O` �ķ
r�gI���fJ�R�V�)3���XNP��d(|����!-��@�|����>����[D�u��D��n��g�����B*?kBqo!���3��zO��|�Yǣ�������C�Ƌ�V[���1����.��Χ0���7�ʏ����d�z��Q�:h��[����,��j���E��l�n�?`�c�	���fG��L��|��bS� ��*�R]����`�V^�����SA*~K�o���Ϋ�dx���<��E��Ev�	&�qc��IOn��X���JA�I��sU���'�W��<`c+8�0*�rL�+������x�&w7�
xY��p����/����}����	C����U���5��5c�8�$��Ϫ�v�����.-�o�_�j��^��遽�-j<F4T�L�M\9����R�,1�\'�>'ݥ�?.,�]�F"7�k	}�Yg��cf֔#�k�p��]O�V��*5���)~�"�:��b>$��3����t�d��#����9��V�f.�өP���VO՞Np6��8��(Kjt���ˊ�܁��oԴ�	����|�;A��|�.؞�3�߱�׊�O����Ot����T��aެf�vl�P�0�y��7L/H4�e`\�R(���v�[E�L�[�`6��b����b�7�=�TX��t����Z2R]'�t��ba��	H��tY^�ߑ��*+ޏm��H�F�x
2CP���҅Ƨ%y4Q�%��)'X~3��C�#�`P\@ka��U�sp���oW��n|q�7�3��&�y�R���ۃK
��ΧB+���9}=��u}��/�Yڱ7�2�y������@a���P�u8Z�R��RȜ�KS�\+#0j��`vb�H3���&�jyj�{�=��NR)��v �s�& ����G.�9��7u�R�� ��,LE}@���
H+���jSj��]�W�{��ӟ�8�j����b>��)E������
BD���=���pL���W\����e���Z\)5�R�tq�{R�8�x3;���8x�M��a�&5����& �o�+9�7£�!���ͥ�|A���-��or���ܗ-=5g�4|Z��M�*h�~��I��	����P�������X�/u�W���N{6�8b�z&�Y��I��2�iM�L[5���d�&i��"�>)�
ET�l�.��L?��/!4��nJ�H���3$�}��`B�(��ˋ����� D��9LB����րD�r��g��떦�Nc�Ҍ�n=Q>�&cw���T�t��u	�*��wi޵l�ݺW�ǌ��v����9��p���|:8�$ő=�Y��]v_��8��[k0P^PRJ�n������t(�gv���};�x��$�o3��	�x�Lٟ|M�w�1も��
����H�p��fP+��-dtm���r������*��g6��E!��{ �l� �Uc-	M��7Ra�C��V@�>}�
��Q�0�Bq����Y�灍:�G=�K���7	�$�P���m���G���Ss���iwg����?�U�ޭL��ڄO����A�r�`�~��J�� �r��.9-{5���4�_���3��r�5<zjJ��PǴRg���S"2\�4\b��"fx�������1�$VhZ�ld��;%l�^]Sf5�����u�=��n('��4�i�$Ԋ4G�9b}
�mG�l�����!��"I2�>��~F�
�u�Ǵ8 ���\��HDy�C�f��O~�ƤMe�e�<����>��t��p'���y��\%0�K.��(�Gu�ě��0nD�a�|�%'\Q���i���R\[P�/E������O�\(��^��J���%�������sJ���;	��c�c֗�sx�lQk#'z
�ϙ�2HR��B�ma�S)jI�����8�ج���}W�/��f:IS+�nkv���IX�A,������Ҧ[��N&P�#ZW
�h�{7�~z)(z�bw��]/D��5��h�j���I<���I�
r��1��O;��d��=��C�PjX��E䀬0�ت' ����I�]{gt��pE5Α�G$^Ǣ�#,�tU��4h��V�r�������灪@�o����=�imv��M�ګ;�i\p B:��@�l����^�as}�ab��qHN
�;��ط
|��t����MVq�#�)�E*�K1�������=���7O�2󯉐��X�2�^��x3@�6�1d9�I�����t6���&�����G�� =I����^p΍P�����b�,f�6�$@�9n?�Ѣ�p�B~3�Su�jy
P?R�ɢ�ݙ"���A�)�)j�q�4���_/�فڷ*P�{W�KD�M�Z��h��*���� 7�v�p�l����Z�t�Ԅ�WH��M��W#n���I���L��ɨ��O@���Kr��Ǟ��0���^�Wq4�Oy|ޣ�SH��^p�Î����d�IS�w�E��<_�Kږ�t�&!�v~��x;+g��y�%\�_!�n>��QX�8�ú������� �\�NS�A�o�����J���v�(���u�v�r���Xn��÷.:�\<�ܣ������rI�;h�ª�a��E;2ȘS�:��
'?\��`�հjF��
���Pŋ�{ɠ�Pߊ)3#�" � �f0R{��:G��]Z�2�2�
��A����$|��4�
�R�K�T�{q/��*�PT���p*y�/�5vJ&���~�^�z�b̻��vV�t�Q|/�w�S��8nw40�VD�O �.��AV�A&�5i�/w�`+���(2S�fB_#-k���;��9�rx���,l�b��>���	���-%��-���L֍�X��W���4�j
� ύ�0Y�X>�O1�'�p����+GZܨ� R���b��NUL�am�K�4#W����E�ϟMBc�{�$��rq��F�P�Yv��t��ޯm;S��Ƶ�b&[�F���� �f�9�ͱS�lwӰ���T�+1ͦ�5>zU#���CH�eUA�X}��1����40�mDEpҷx��\�)W���`��	W����|���i]Y�P�Nه�����I\Z�M�j9��"vF�;{�!�m�Ro0a�|�7���7
���6:j6�/S��*/&�c���q��Lz���%D��Q�~���+�'�JLdK���n2*�HMQ���΄����i�d��n��cT;�6�[=�$��!>��������fPAC,����J�T8,���5���,����7�8jå,sE����������+4��߶�M��6��(�2�)g�#ǃi�;X�`�XI�?����߭�Z5 ��$$�` @���4��t3��ҿm)���8����Ib�ssaG�1N#������������?���/+���G�j��H�����qZ[�R>���d
K
�?��:_ġ2��ѭD�P9���OV�K���N�H{���~s�2�������+�j���-��=B\y/�.=LK������wX����[N�搳�W�DA�4�]���iL�k�ڠ�;.�����^*�{�L#�{����N�W�_�"���O�ڣUP/j;J~C:s����/NXf�+�Ĩ�r�:*%��B۫�}�	�K�h�oVh7��|t�`����f`Є�^3-lo+.��/�1� #�6E�j\;��|�j��c1ը�
��\�����F_�k=�%7t�/#:�M͘.����u=tO^W��)���r��h��'_.�����L�2;�u��wA���	��#�U|��RP�'͟�d\ܕ?Kd�2'J\*�cpݨJ�{ɿ�<+?.���f������^W��dz����!�4�	s�|�L�#�
of�������IB���21mlKc0�(�|��y)�����a�=1S��/�~
�����z�dW������w�X���	�y����Ij�JGȐe�'g�6�,F�G���0@�MK�6�(��	�ue6��v� ;�٢y��+������]�bp�����~G�^������j�L�k+~���O=����P����7�k��h�QB�FǞ����b���7mۄ���uߚi�?����kUK&q�tޡ&��*i�4�ײ��(�����{��յ�N��A�c5�����Y*>��(��U0�ʯ%��k4;omT+��|b^��]�c���D�y���o�Vu��qݻ�XV��?�$���{U'�Z�mTEG��f�K�����A�����+x_����'Y�8g8��A��*��.���R�2�Â��&��A�KƟ�1�LS����̬'��*�'��5V�u�%�dK��^�3g�|�"��7�XI�Rs51���u�糀����o$ɕ�Ɂ�q��$�v=|��?N��YL�_�^(�X~�T=��53L��M�.���.<� �:r~/�2!;�+f�0k��`�Vɓ+j	[�� �
ݣ/7�kBy��}݇ˡ*x'�1!��MW.ʗ�;���^96���<?��1����B:�:���u�5sϫCqP�^�Q�?�Ҡ�ʍ=Qij�
D�X�2�����e�q �����X��I��s�.�_#�< �G'$ܧ깡��i�PKJx�0�J9`�g\Qʗ0�U5���g�� {]_MO������~5us��{��1"�*�7(iaѩ�'��A��i��SYڝ�\J�A�4Y,�RԬ�򄕓|�����(˟}A;(���;a��3�_%Z��5��M���b��B"!;w�L3� �a�]4��な��q��w,2���q6��Ғf��E�tdtb���g��R�(�M�F鶄�$�'B��@b�i�}^��@§0&v��zg��66�B%��fi�l�;z��2B���V[K�b���_*�����9��Z���IU��ʇJ�c~����-_@T?�$����Lb��������@	I�9��띇�F��"=.�i^��[�N���'��gr^f=��i��۰��meUk�BY`Z����dU��t��֬�$W��j��
�V��R�p`��̾�m����Q��i-]�K��Z�p�#	˼��%gs�Is�dE�W6k�@����Y�w�ُΎ5kx��6�D�
�'�l纥un�P璀d��${�̃���_9@[O��Yh��r\&!�u�nt�.{����Qg���D9*���ƒ٧i��=�O1�����|��*GLJ3Dr��\%�o�@����x�6u�C0�(l!�I�#���Z�X.�c�(8�����6-��w���/�&�ޕ�+{�>D�^��� Q6@8���Z�=`�G`Igq����Q�_�����L�Ld�u���vכ��?���4���f����2
R��|��s}�7����)L�d�l����l�����ڲ�ͽ�܄x�%�S���<�Ο��{=+���Ă���!0sg�����e�`k��N���O8���;��Z=��hݱ}���׿j��یLM �[.�,2!-��eT4Fu�*+W'6��-����t�;;�"�~�_+j��ݽ'��;��ǟ�a��	��ջPG�21�[J '̆F{H2��'CowY�'<�f}�)( ��k&���h��a�X;���BI�cT�#�����B��}خ��2t���c�����h�c��Y1�űr������d��ͦ+)�.���Z��_#�vF^�4�4�4gdB?�yˁ7�C(=*~�X�L0%�� [�e�~��:T쌹���..R�T�K�ۓ�Z|��R=���{T����5i�W�>P�����^В�h!h�F)�U"q6�lC�c�@��j��
��n�i,sr~~(ȑyW=ҙE����#��.��]��dN?�&�s�B�����<���@K0�T|b�(r�D1oy�J����'���K���1�X�h�
,N �Prg ^ܲ�-�m��LQ����Ie܀�b�#v���:��~��]�6G���.���}�o�1��a8	4ր�� _��L�qiis�x:s����*�c�N���OH;+�A��k��n�rwy���a�:��}j杞�&S���5X#�W����B���80��kM��/���K�q��ձ�Yr��W����0<�
���{�-�gt�1��{�?���m�4��*��jݢz��w�|��"���#�/�b�+�Ӻ��]��?�	���s�z�I���[VB�a��1yH�C,�~zlyn��.�Z$*P� q\;�ޙΦ���Gv���	R�IV�)��X~�Mex������ ^�Sy��NKJ��3��C��Z組���!�	Ҵy�*n�]-\���7n��"{���ZȥH���xD-U�RI��j_�����7W��`+�"��
�+�H2L���X�d�R�?�9�����y-�����К�O�6Ӈ귺��P�"[`�l�k8]�[e����Y���RɈ�p!yFV]��+B`�z���:E����=G�]�����I��ndG�(��R�H��~�z2��'��t�R�q.%�����>�nv
�&{j�y���ɣ+9M�@pS�VQ�o�d*�׶{�������ɱ�Y�l4��g��(��;����y�0^��jv�X��]����������۫K"�+ob�)o- ��n:�f-���������7���a����?A�kWzT!��nP�.�"�H*q(mvEo2���
��%a���ɦ�VeE���j̠�����SkSd�kdsy��2�M��� ڝ�����I�ئG2�Q�V�[�A�����J:����i���&�t�<��̺{>b4�����n��U�K�o0�8_N1�w�B*��,�l=W�4fӗ��\W3�O���:#�#���M����;��%�x��Oc�%>1O<��[��@�t;��PX�ͅ��P>�����Z�+Y�m���$�1L��f�yK��E(�N�IH���Y-��[:2omV�O[��8K �RD�J�Vb�o����k}�A�������(Q}����K�5-2�L�j���GW����ӑh�U���b'�ah���yg�NK�IH����,��<����ͭ~H�tGЃ�y���R�K�C�c4A�Ol���'馾�ǰ<aL-���{�46�(�C��!�o$�0)��\ �P����Q ~jds~�SL���	�W{A�	��U�#4:��;�
͆_i�zN	kF����4�F=X�cw��^埵Z�s�;ʸ�k���e5E��<�Z+�o�׏�Y���rS݁m+AɂIW|=V���:`*5� ê� tRX��O��6��$�d����Q��� 
��-Dh"~�����~Lw���0����]8��H٦���H&�z��(�����5;(�t��K����VZ(�f0ò\�_5��u36HA�Z�S�hz�r^.�� Hm19J_LJ�]���!"��_1�s:�d�[~��V6��>��~�� �+���I�Q��s��P0�T��ØWmaJF�_9Ix��o�������qҘ�7nZ�P�������{�|�"�uu�2�7�0�qw2�Et��T7�5���[F6�YC3�7�b�0��PQ�شi����͍Yҿ<gz:���N �Cϰ4�E�P�Xs2w����ů�������5�#ғ��A�����ӑ��E���z���K�Щ�z�Go}�+#��&f‱C��h��@m�lp�m�PFE�*tvHh�4����gk���JO��zÂ�)�6>�a�?t��8�T?i%~.���i����^��)���� ���K���Ge���3�*~�#
�������ՠ`��*|(��چp��KiB(�/���f�@7��9YLw����]/��X���%��`���Y����<qD�*��A�T��jt�@�w���r�W�1q��=���hT���%-�j`��us����N�bg�O!�&�J=��}j�˔��#<�_�4$���8�kob�������:W�W>�u `�{�:�q�D�9�F������֬D&�4-ć��;�?�N��F�q Ԏ /%#��cw��_��i��\�@�4�(3�>%^#�.�+�%FF��y���M5\�&�-tԖwD��Wp����k�I�T�������)�������CN �*�� ���5(i%r���ut�Q �o�,0��ڑȧ^4 ���1A��Pɮ�z��]仏���+�[sI�=��Z�{�%<ש"�~$&Έ�-����z��Ts(�B}_ ʜ���1�O�9$�s;���E�������<�4A؉�����X�`E�\���c��� &F��4vJ��`7j��Y�e��h�U`��ʌ�E��/"IK\�RV�s���[���C�`�\�o�V@mf4J �֩t�qg�a����h=���K��n)�У���("�~�(�/I��mv�����D�ѐ�,�#'GmJ�H-|W�uCvrSX�@�<���A	��&�c����-�,����S���!M�0hI�7�g+������x�H신L*���?az�v�4IRU`"P���[β�v��e�.����
E�Z�)����-$�ɉȳ�D`�o�CJR·{�+�}R�#�ĵ�
�k�;7Z�ݧa=�L���q�����N}Ri�b1c"_gT8X"�ϙ*Vv3�������3�d���쨉�������m�����9`5s�|L$O�Y��0���!��%�ۦ�Im?�ɹ���p�PT�$~w���J&�'1�%���}��O/xX��/5�A\*d�Gq��v���1�Q�_��]�_�'<��G�ۇ:~�7O7�����vI�G��\����C?x�!?��]U���X����7ª�Q��@jR�<��-��H��*:��ȳ=�&O5�·��V���>�뾕+k�@����Re��6N�Fv+����ۋ��1�{�9���#�H��ވ?�i��1�՗O�i����2�� R�����K����92���4�����W���2��"9h�K��#LT�W��0WKq�ǘ�3�F?��DF(7��Fu�dT�tj���y�z���uf�T�e�shzZ��"���V#;x5���F�-��߿Z���ٿ*��ME3��᧬r6��Ϳ9�'��B9?#3ȿ���8 �����L�"#�у�{&gZ!�[��챍}(�=���#?��rW�߽jʻDǄ�;J�lg���<��w5D\�ʖ"(d76�=�?���TkU���ݛ��}L\��K��4-'�|&����9�&���*|��q��5�`�p��eo�6kn?b�U�t3�p]j�d�>qJ�R��]�7�I�ԓEs�Yr��eR	�Q0:���d�U}�p�5��-#tNC�ѩ$�?�/��N�t;�2x���MG0�@����./��� �
ȟ��D	|�9��B�^WZ�K�3i�q�����M�, O�0�Ю
˥�ױ�o�DhE��M�Ӷ�#�Ơa�w�������E����r<�R��C{��K���Rg�䥮ʬ2p�Am�R�@ ����IX�*���0��t��-	��dX`���V�d�ǔoDX�]�VM+�Cְ5M�����5Ӵ���]�5�kJ��E��v<;$v�d��0�T:b�9C��k�}!�;�Ȇ����'p+��k�$������3�2�%	U0�v!J�-��+���@�4K�n��a��<%�!U�3���-fA	b�����GS%>(z��>~F�<�k2�O�P���|��-c6��C�������Ҍ>��`n�uP<p����hNz$�~ˑ���Ҟ!='��p��f��2.�!b����h�Y���m�G�ގDy!���x�6�����H���u��xu��ULq���_]D� Z�X�8ި�6Եt3��/�kWh����Q����;kN��S:� �U�aޝ��#��bI��%�L��=>����v��~̍�~ș<H+P?�K&W@�����2��M�}o-a��d�i�Vd��	Tx�2�>VJ��G<T�K] �����͜��>�\�(v��3:v¥���c��wo����n��f��l5
loD���I�`H�:Akm��)O��:<�����m�х��T=��q}��!��;�][1���S�ퟞ�sE�0>�� ��G`�U�y��VX�9(�s9 �4���o+z!�.�(H��y��;N�B )*H�^��I�B�-�cT��Ha��㹖��v�
��Ȥw"��m���[�a|q �R��iZ����w�̒�W ufV���C@|�T[ė��ޫ���˭!ݞ�．��_� ��Y� &�X��I?gbw�7�K�ΨZ�H�	v�x��Ϝ*��R= ��E~��׻		�4ѝvMgx��4^��]6!bS� �,��TBn	ᗯ�6%EX��[�#(K��],AI>] ���.)����_zn)�>M��P2a(�@6����B�&���Ct��
�%�Rh�	���N5�Q�*{�H�6�O�5��:Dq��7�e������:�R���m�tx^��gz˵�b.{]�C�Q���L��c���[=����0�)�>N������B�ѯ���/<��S�Ͼe?a�����,^��K9����9�\�`�ϐ�6��ag[�;���2�V)o��9`߹R�wWsw3�q��2;��9<�Y����fs��3�D�/�c���
 3~gU��*@Mx�'J������jf(��i��A����}E����dW�4'�6�Z7����B2`�[R2f�N�u���I���!z�^�1���&㞨p�����c5Z`1�~���k�-��VS^�����Q�	����$�x���)zq��Ɩ���7��PԌW	��-�`v�^�e��~��BT�yo���Q'�d�H	|P�J!}l0E4M��&�U��T
��gs�sRY5��I�����(�*�/t|�op�g����~�j]�B��,�XU�n�!X������l1,Tsx���\��������݅��	��x� H��������Ҷ�h�?%t#��/޿�D�lҧ�)(^�?�<
3z��\�q)D�Tp�4�k�;	݅��y���e��ak�k|�{�i�L	�Qz����g���0�������X7@�Q���;c�?Iq���KV,x%�B��}�=����Wn.������5�U(/$Y�����gP��X�HY�~�G�������Wd(Z���J���0'���E�f8diE+:	v�6��Y���p��9]�eN$Nޅ4���V{�4�.Դx�Rࡏ^��S�I�K�d��=�R�N)h�,,�Ao�k���߹�g���}H�˅_1��$
ʟ�ۚ����>���6u����!Qb`-٧�I�z�K;�D�J�I ǆ*�2|���f�Qw�� c`#x����;��W���sּ�s�P���[yT�Il	z��ec��m��ʛ���<���G�&(��RkL�Y+��=�
s��%�MU�kӯg{���]P��bX{����d���t���n����ĻZab[��PlM��Jʲ��}Q�(���>ZY�E]�r)& ���L��WKvo䷞!H�Ϧ�Ҟ�Q%��"ږ�r�.?�yG�=�o_��}AN�H�q�����Lm�^�gC��0�I��q�@��ˍ��R�T@����u(�:���`*s�&5��dbt��� ����%�q�6�.<37H���)Ⱥ6�9K��5
@(�@!�%~9���v�;;�vY� ��ݕ�o��Q$�nS��pƎ�g��n�ּ�]7���6�0(�#��cph��FRA!:����a�|	>� nȜ�k�S��U�������Y�{>��N��N%����{u4c���� �<.� �W��c׉�D
 ��oHF'��|�������3��O����{T���C
�m�i��6�3i��Zd�>���r����9�5���.
-:ѤD�a���1R��e��R�:v��-��v�+�Ɠ�۱sl(�Y)��dO���a8��8�Q��6+�Ъ`�8�ؕZ�c�$f��4���YF�RW�Qe�P�ʜ���v-mn?�Z� R �>�_�L�d�C!8��lV���jT_I�7��L�?^��#GlpBb����%�闷`��ɬ�`2s�5K�f�$�(��H�T�E�Sgζ���ζUg���uCˆ=��/S�a�r� @�|湪�YX_��Ƈ�m�C���Ծ��~��shx�8q��^�t��@�I��7M��]8�X���Rx�v��s���V:M��$�����8"'(���m-���x�V�a�T/����B��6��daR9G���E�n|��fH�/@�c��S�}18`�W��@��]"2~G%0l[Ҧ�1)m����Dx}������x��ʯ��fs�;�Yy57S}e�����妵^�����#q��G~��%��X��ӈ@��Yt6`�I}jO�f�#]{),��5VI� � �,���~~#>,�cZo�����f����y_�x`t�W�ew��:.ȡ��5?b3��f(D��7K�hB�h�?FT@Q`L�8�_(�|�O����H��9 -�t ڰ0`1zBn�I:��2=�덒Sq�����|��gRnWF�u�[�A	���I���DHY�U�u!�Ey�w���u�i��6R�t�Wb���f+�187+�^>1O@f�Ɛ���7N�ӵ�ap{L�$!r��aB���J��x$����P�@��@ܖ�O_o��������]�;�b�N?�jx�\Db&xl Iͫ;�R�[Q�hO�༴��dZ|Gx XCK� 7*⚔���K�l�, �ܛ��@!�J��yL9���$A֌����CN.���׹��?4�\5�:m�G�$�	���N���X�1�G������_q���j&��$�yu����p.��E�6\�^�Ƹ�'O������w�
�YM����QCD����E'�(��^�
5qN�^']�lUp��SE"�'�����]����=�dgW9�^l[#�0$@�^bW��rt�RA;U�٩V���~C�nY᜿u�
��A�T�ܠq��7����w~e��z-�?�h!;Lh�V��c�ʮ�1D00�v�g�������(OW�жN��G&y���J���$�o�d����&����U?&$�g[�kl��^P�"&��%�t�~\a�YF�3h���Ψ�Զa[*�j��|��^(�
�7
��h%X�fk�#o����Qћ7F�58�Ƅ������������='C�
�����d<�R;��hH^�f
ƦE�� ����bE!^/^��̝w^�)ޓoy��(���H�:���P��@�~\���[���lG�&|��=��9�OU⋅b��it�[�rY���	U&�t��N=r��mnY�{�U�/��-���!���E=:|�B(���;=��o�����m�I�87�Ó�:r�����S�Տ�M�v+Bprl'���&4��.:�*|t�0�Nv��T��+wI"y2�T~ǈ�i�6S�rL?��"�;)���K�w��`m�d=�g&Wy�}�ϡ���ɉ��#u ��Q����Fی�?��럗g��˩��|ػ�h[�Ǵ���Q\�;3�"D�P�x��~�a�2���"�	���
����<4��1Y�e�<�hu~�衋�;?����di��Ow68E�n�9� $��|��Ta��c�<�]��T��4C��;N�W( %I���<�Y��U���&�G�T��>�$.w�i4�(/����G��F�f���WƋ����BP�#A�*���y@,n0Y�����zc����Ëb�g�2�>��?��O׈�O:&��K4�O��X������OE�ҭ�e��,��"㒒n���W�!?�U�1�k����u$�D�1�x�4��:v�T2�w���J�n`!,���Y��t��|x7�1;w??�<Q ����{II�k������E����Y���i��e�wB`/�^`��Z g���{���C��L$��,�2���O���ᰌ���e�.��;�=7�P�'[$؏և��En���S�*s[%�Vez��[C7O e�^R�r�0���N�DYH��I.��G�Qv���|���dr��3��`��PB�Eh��`<G�H�딽���zX:�O�\*=_�����V/���-5���������?δcRb�����JC�<�$����U$�yoΪ=��<�?���Eܻ�5,�煻�~���J��#Η�\��'���'���zy;Ն��?id�5���{ߡ?�7�� �5g������;h�2���S!)\�e�����ص;?���7�>vu .r�?�$����9������Q����bB��[�{)��P�m\��j�����F�Y*A�Gb�H�H�ާ�5S&5�Kd4����PW�b����`�g��V��]MƋH!wT��%����o�J�A��(�C�K���O_����|�C��I�7�k�v-�Q�^9�n��%�jӟe�����S�I@��Cc��>]�O��K  �(���@|��f��\:�Z��������p�K��h�?�K�L;�5 �KɆp���2�Ξ�}V3�G��<�������{�!����6s}M���%U�=�I��'S�A1��B���Esȣ�������Y�ֽoO��6÷�6C֝{�.k���6��`� �l��㌗��;�wī���4ә()���`��� ��n+��N[z�6�).hb�`cC[	"�g�3ś,��|C���ҹ�*�mJtXZhYa~3%7�4��c�r��@~�tE���a�yӥ�Ы��� 6*1-gN��DU�]��&��1��j/k]�D:��ʻ���Ϊto!�a� 	< �����V�uq� n1���DQ!��F��!l�ڛ�����բ���3l�B@�Ȍ�*�v㚦�(�B�&���*�t���W�;�P�~�xl����L<�1g�N�s�٨���Z�=����mJ��mp�ɛ9��y�%ׇI����ģ�Mz�o̧g�����l���|���M�6��1K��I֍�C¶3���1jp��ŒYI߁�w��v�N<�x�Š���[�Kf�8F���*�x�u��Ry�e�����cp�۰+�MUB�M�#$�K}5�w�q�R�bPé���6)�����F8+��^�~�	"f6�P&HC?����-k�J�վ������%�-msO��6k�&W���t���(n��o}Tapa�o���  �OOfa"��Rz�)FTB����Np�=�L���G�Jy�
���b-*G'�K��9��"E(@[���z)�� ����Y:%o"���{k�?�D�w-��J�J��]�F�������}�e't4s����ס^���GW�:7����oĪ蟩]���T����˹�{��@%	d�D����q��)���������l,7Ȩ��B~]�K�l�2d��!pGU~�ۋ�l���"Cs/���͖�;'ƚIz�~UkY�[T/+��a$�]3����:+�{�(�C�fh7��Z���С��6���C&�G�x�0��٨��ul�V鳊����E�?꤄���6��p��J�ǿ:��Pd�k�6Ti���2�fT�7�1�:�V@֝porF[\�f�����uV���pL\��h�Z�zz&I��*��jG��Vkh��.�w�m�)�$3����H�(�xN���� }<�d��+�����<�w�R`L�&i[l�-��'�r��J�(��A;&J�o4Ho�It<)	�o�y����?g������p�.u��$����vv�H��m�g���R;�������z/|v��i��b�����#����PP�"�[%�o0P���D� Ժy� ���8�C]\���"����2@WtȀ=� �[}�d��]�W�¦��|z����V��3��`1�Y��Z_�*@�K�zM�+��>�J�ġU������,mW��>�j2��NЃ��_����u�Or����$�u��cffb3�S�Y��(m,u�iQ�TP.4����p��KT��Ί-[����ڻ�Aϩ����;����u2�ˋ�K	�`�$�KQ�eL�e����sW��ZYp06�o���KaCH۷fI�b���'I�^[���y�;^*��`Ⅎ?�n������}<�����	��ͳ!5����0Ei&� =�b�j'!Zvi�)DX�]�-u,�E_=:�	�E�E!Y�Id�bx+b�I�(p�8�RM{:I^��?�k�����D&��2��ק�������.�(	7[�;=�Z�!�!$|����!��\�L���`f�R�
/$vWegl?�W�KA+�����k�G���x?A]�2�R�h�nV|µ(B�UfJ1#�)��(�R��h�M���[J���]��j�2N��lR�r3iC�n�����f�e�$��0��#SD���X^���	ɍ���aEfk:�a6+d�<���^H�/�x�,[�#T`;���%zƞܯ��i6p�؇�5��ϑk٨Po?�Ԕ)����x��`�ar�oa�S��~\��5�[ ��z�􎿿�Q1v�$[����C�C%hL�9�^b�~���7U��tm����,�ץ
T2���Z�!'�c�w�ٯ�j��яe�`��Bj���y�]П@�aK{�fʻ�Wŷ�����^]O�9����ᏺ�lO%�&L��3���7����Jf�f����)�o���� ^_�w���C�7δ��'�߽�3�uNFm�7bI��|���r�g��o���XHG޸��zuK`�理Q��FW�T®�pH�� �w�� �+�%dn�"*R�M�Dξ%���R/-,�d��YX����;}�!"s���e}����Ɍ�q��){@h�F6��2e�܃�_x�zZ�G���}�m}�̝�m�}����Ŝ=( �L�,��<��CR�'mj�i���gw����cUfVO��$���$>Ui>�^>{�V��,!L��<��KU�
/�b5��T!S婊����"�I��@.ڥ�̒��:X�S��[	P��Gf��=6���2��U��q�A5��V/	�c+�b:���/�Z�+�.Uؕ���!m�hSU���ʆ�5��c���[�>$yh��e���J��`R�uO�j��Z��h�rd��UkAr�Si��K('���}�zHfR]��G�S�)�/�Mv���a���1d�O� ;)Ϯ��"�N�1��LmPK�o(�v��K
? '�}��eS��@���u����4qK�^X��� �< 񅭬�pQ���,9h��&�&�5e æ��i^ɻ�]��M]��=���Ť�ġiKյ
�� ��2����A����
�K	.��~�*[uPX��^�� �(��=?.�C��)�Ⓢo��cn/pF���>@��a_�W�w戆�����v��R�A݋��Zx��w],%Tѐ:|���#���2�|`�Y[��L�-5��ƪf �S�Cq�a� �ɘ���7�������?��x`
�RgØ��{���
�~�������i�h�=���+YF($đ=Sw��G�u�B�0�}s��jP�X�P������gd`�D*�!�r#�o�ý�^W��~ Q�&��||B�Q/�����膓R��gRl.�8q��C��*�C�
@��fup�#�?�:5�3��i/��,c�A�	w^V�Ǔy�Xx���ZX0{;�Q� ��]S�Dt�f
i$r#�<ӥ�m�v�!�|��=@��V����K�2�%�{����H���1P��z��Պ�/�����ı�������$.��!�x�n[�c�R��}����0��9MI���ٛuFd���d��x��, �Sѷ.��~rJ�*=�X~6�'���'@"Ps�r9>�F%�fӈ�4�f6r���Ӷ5J8
�{��&�{?�h�t$�\�"u���(1�p�4k�}�t�ڹ�}U�(zK�*(M;'݇�=�gZ]����a<� �;�-�-���	QI�_9�5� �����T��/�	+=����,�q�<@�-Xԣ�JX�c;�zU�;lK��	�dr���<��ڗU�| ��IQ�QNyЊ�\�mu��qg�؏�I���S���ʢh�M]����T�`@��e4K��DQ�8�>ݐ��W�&>-Y�wQ>��o~ϸ��)`H*�ř6^gW���V8g��/DͿ��2b7��jiDH#��}�mXY�RQc]�U�'�H�����3���p�Q��w��#���Ϸ�50G	��m�W�7��=]M��Rb�_�W�O��c�Cv�O�[��It�����%�U�E�qͨ���b�|���x2N��D��_��ܢ�	��,���J]�� ͝�T��������HnS��8�$w������:����J����2�}8ċ�ǋ��r�S\Mde���a;����2���b-̊�k�ą����#j���Z�W�<23Y3��1�5��1�^�tSdzΆ:��M������@�C'Q���8�YgV0�Nɢ������d�R��RV�)0�qڦOZ��4!2�Z��0��� ����l%��ޙ�L�<�����$�z�k���:�R��Yg���Q֥�P��qiG2 ��)��8��g��cdt��^ə��HВ1�f�	G'�_�HJ=&�GO$8�N�A�9f$�B�6�uH���Y\�im=Oq�vۋx�O����*}��v����}�>���wo 'q���~�ӊ.�tB��8�si���}�Ű�#YY5��Z���]��WGBy��,G��S����ʝ� �4�~��?+��r��Z��?ڙ��� ����<c�q�`\vVB��~����go�e�t��d<]
 C'[�ĕ��e������'�/��Yf7d�+{��L��bj]��.��zUҍuԑ��D��e��V\�[��e!�����z]M�sq��l�:DM)J1���(gQc�U��LM��A"��n��zD;-�r>��{��u˂�E'b)P	P��F�Nulj�b�뤝�\�F��x�"{�΀��i�N��T���������|iL�jr�fG�M���̇_u7�4 8��8���ˋ/q���K�J_{��n�T��	BW��P���$�P:d��I�js�ϖp�Y���S ���x��hY���~=4ӲH�N�����H\re�NR�&㊼�ɳ��(�Ux:FC����!��u+�tW�_���y�ۉ�_]��eVtg�C�TF���;�	�g]QX�(�g�����ȻX�kߔ����P�y\H(_��u	����KF��P�bْ�qv��?8�X�\�Q.��5S�_�'b�C�m�	��}�KF<Ԅ�a��+�8ӗ�7@�v��[k�akRm|��b�?��:m~�����1����ş8���&)D�g�_;��g���e����ߑ��F��f�^�Ϥ#���3�7�������� G�e�&��RJ�=du���kl���$� O~ �rΏ���z�XQF3(�{	U���4�1�%u�쨾�0�17*�xڱl@��������3�ܤ�3��=g� ~t�s��vyOEr%�AC��H2��T톁3sy�¸�,:�pE#�lj�m�%�z��Pu_!$n�iҴ��#Y�P"�p�l'v���߮�Z�,EZ���}��t�F�Η $5
q���Q�mB��=�a<=\�1�L��l�M�_S���^F�'K:�.w��g�;5���ae8��)�4W뢖�G�ջn�4&�Q���q%��bͣ�`_E�Ʋ�����Q�BIU�H#�i�Kh�U��������b�h��O�6�.�{����晩��Q�Y	�+oL�N 8-np��	�^
� Kޙ$2���;;������C�ꀐ��ι���8Pv*}�
���K�X�N8��o��F�qS���F�i�Fgq���(�-"1x��T�{$Xuc����2��N�a�j�*<A����4|�s�	K�r{���Tn(� �:E�_ͤɡ���ư1��p�_!Z�uL$�ڒ�*w`9��	S� �[d���#@]ҡj^��prK��nV���
d�>Cǟc�\�i�B�G�b�����h�&�q����j��4�����J.i�( ���l�O�mR=kߠ��^�PP�5h�S)m�m(�ĔQ��$)vaex��ꐿ���S'畴�b���Oz�+�$��{����w8�*�(���r���٩߇�ȫ}c<A�	h��~
Iss ,+ﮟ���Q�˵y�;*.���4R�$�C���2�Y%E�+���r�{�٢k���<ql�R����`}sN�ܽ��0�c_�1(�C��7����k�����Ccz@���ȹ�0��4s���2�Ѕ��������K�
x�j�"�Mۂ��l-���j$�>S�K�5��������֎�&q��q��	:�gWUh��z͐��[�I"sN��}��=�4ƾ�?�.��V�sشƢ~�jƸ��tR�U�����v�{Z�[X�.�<�/�8(1)�Qܢ�CʜV�p:n޳��l�ŭY�{� �EF�@b�q ���Ք��aNs�ɧ�t�"5ӽ��$?����ꁈ��~cuQR�J%�U�'IqKP�8�5̧ËԨn�����z��u���}*�8r��_�F`���Q�k&X1x�{I��}3/�߽�F`�� ̃�;C���R�e��i7����XA
�'B(E��������a
�A�Z����M(0�<����`w����"�j_�m��ߍ�c]�a�<,pYڎE��Fh�̃���3mZM�u����e��:�G�P*4O�؜��O�ָ�-n�mj�H�at�E�H��o��2�b��?\/+�=]���ۣZ���A�� IC�� Č5�i�c�:1��'��n;*��J�� ���p�L7��(7�\�����u	'CwmY���	BL~��33�:z0h������"��R0*�#����h�����jk��0И�B%ϭ;�C��p�������	�����Wɧ�:q��7,m�֊ɵ���;3X��O�'%���I��Hy�G�*�cm��LP�'l�)_u���"��{����9��M$!h=���֣�>?e��)<� �Z�TZ��qō�#�"*��n][?7Y�Pղ�V�Q�uND����z�EPD'E�u����m�k�Հv��5���5���Y��R�9��vr��.Y��y�+��"�O@�bGB��Y����^����Zl�%wz��P��«���F����-�g`�̈s����w\Y��W?��p��fQ��R��:��uM!�{'�e���v/2W�|eK'QB泼��2���b}w{�	޸��%�F̀@��P�[���b�����.|��CRB�k��[ �I�s����P��~���#1�g&��L
�!�� ƕ#~f<�1� �ahO:a�V y1�wj�)��A��]�#��c�"6#�+1���:�E�J�u�Z�A �dr�<a-�[�Qjn��%;Vtq�͉o����)�RGRC��OS��W�'V�\? ��� ��)
Vj��nxId�zU�+>9�:�-�������%,�t�$����ͭ��y�pp�"��r����l8��|�N��v���Ma�E��/���m��4�@,�3�y�����7d�]Kp�l|`@����K83@�VcH$�=G��T\]J�]<��P���_�e��6ʰ*�_�ߌ���퓾d�At�\��A��Y�=�t�Ү����VO��c���vL����i�cF�@�M�#�Y�5��A��P�{(ֱ�2ٱ�wq�rg� j�n��+�*Bל��?�
8��k))Ϻoy�#�A Lh�<3�OK�/�8B�#7A�K���y�+���ȹ�S��%�<�B&n�.�t2:�i���{�m�o RF�@�|^R4�$�� �V/�z���*�s����}����f���(��ջ�ې����{���Z{�t^��_��i'KkU�K��ڧ���PL���^��;��=�/�T�08�6�����+5����l������/�a�$����6�4�s�1g�-wۀU�~�����p�gRSn�;�!DL��z5ɐ
[@��
�_��ieB�y�૵�FKԴ.��	��h��^�a�{Ct�b�z�Ewı(tu�5	�K#���VI�I^o���ů�/��u�@& ŷ�JQ��L��/�����o�T���;���,�E^�."� �����2n���&�a!x�f��y�,]��A�S��Zf0�)CZj�����QRd���'48�ˀm@���\V~�i+iQх��߇�_A����zе���$\I�d0̒�v�U�����8�#�.�~f��C�)5P����{��l��xp����a���o%{��G^
놣�*	����C������dL��J<�����j^&+�PȐ����m`��?��-�3��ܐ��N�p�0V7��΃�{���w�m�X_�W; SH��s��PV#h�9�Q�'�o^����{��
7����f��'PA}��r�{�_p�j/񬞰aMn�}N���l?^�5����,�X�%{�%�����pո�KȌHὝ���NTe��{
��|����K8���PY����H̕���_���W<���I�0o�xA�j��t#��6+u�]	��~�3j�ҭfWP����s�U��$pNT8;�,h��6V����(�x8�<]E�=eɜ�YKeP��ɔP�,JCEлS>"w�K�)���-S���_�c�~?��\�j��\�$�FW�Y������M5Ҽ���Z���r%��lhB��)!�����;s&�H{	G%V�%pQ�ԇ�&x�Uh�@�E����Q�G1ՠ�t��=�J7�����M������ka^v!�����y�f�M;npR����B8I��M�M��nBy,�D�D)t���'���}l����]�z�$:5�Hv��X�c�TW`F�V�{��f��lp�ur�m�Ő�� ����Zr��G�2�̃�$��N��(�:��T����o�5ߑ���oeΰKj�)}�"�ם"�mW����hY�0�;���� ��� ����s��U���m`��98(��W ���ڃc�͝��:o;��_��kK3�R���[�,�}�?�p�����T��8'�	B8���{��QB*��Q��/ezy ��(��/ %�z���EԮ�)�B�E�Iu.c��fÒg�҉����?�d?�ޘ�L��4`���w�,�-l�1��a� %Ȥn�5��7x)\��3�j ��j,�����ԕ��!�bj��8k�+$���r�LG��Gg�;9 ��\�k`�]=*�S�Vܻ+FWs���>���i�څp�MUJg�ϑ;�@�a�/��ȭ��^��yu
��+���⯔_�#b�h#�u����R��q��M����KyXCتz���)5>K�6}�K�h'(y�H	sYmcg�i����C=��L��:i�b�n�Rc����}	E�f�aM�:�p�w<X�`�h%�>��R*f��*B�/����
t�DĂ���̅�!w������������ʥ�|ېH��	�2Y>�Z,�(�/4�G~���cX�\[~"��͟	�rnׯ=���B���`�%t6\��o�G�+�6�,�e������!_��DV�iF�p`)��
���o;5�����o�([:�����Zd�o��g�(9����]�F�.���I�����`>r�=c(q�}��x�����Ŵ� /���
]*mb��L��py!���u��f�� �|�����s(YB�/��:�����"�8�bk��������l��ͯ,�a�wR��!j�n���Xe7|�σ�-��!9�|����#�;n= �����1���"ِz�%�7ރ����^�V�����<��2�$�@Π�R2�{�SG˴\�t����:	3-¢�y�o�i�T @wFX2�����j�?~�}��0��0��2K__�ȑ-�b�ʴ,->zA�����#�����2{�ԮG��E��4���H	�dԭ��~�iC��Rh�s���,�ќR�ժS0��J��3j_����B�����Ku��F��h6����{�� ÷h!O3%:��i�2��U�BF�ب�ѥ̏�uҾ����у���
̰�ܼ4Ҩꌉ_��udQ��b�ߴʎB_� �4�P�Yot���2Q`6P�<e���I)�9u#�c��c7�֞����jE��/���P^Dg|����G�����b�o�A*��]�����V�X4&����?��ֻ���rw��%���fa�P?YͬW# K>���W�[�i5�>��z<����F	6H-G��S{۵�/̪`�߳���V,.@��2��,��
6��󠼥�V���nE�'�5���LE!H�aH�*�l2��<NUP�Y�^4�R���h�Yķ��#����\�I����b�H�e�.��B����d]:�;��$�=��y;�>�\u-�E����V��}d^]Γ�"�ع��rM 9H?�n�)������v+p�~��Ƈ/���T��2�;f�����$W(!/]����B�?zTCp"����;�N*Ir��7�&֒%	A��}� �+�%���gʓ�\\�j̖����Ni�g�7un�	[k=��d�al�G�{��=	��j�@�rF���'_!*�&�cE)��y��k���	�t�|���!��X�E�\� �B�B���C�f��?1�h7ا�b:`!mQ�����%�&���YOuƼ>7��gzwq�l��2-�X�qH��`!$#��U٬�-m���i�̆�}�0�㓫�|j�?f��Tw��"~i&j��y$t��K��1Ҋ�8��t�%
��}*����}�ʴ2ѪH�5��#�ҩ#l�;������Q��Xzd�|�e�����]%Ws��d�z���U���ggrlc�eiO�u��������E�8�q.l�N���xb����unN�N��dQ!�롉�^۱�˸�.����jk���6(�? o��c��zy����FY�Z!�V�R��Q~X�K�H����%(���+��9�f]]�@IY'�B±��1����hFS�"�0M��P��{�z�I���?�>g���`M��C��e{�G�/�>�E�O����qb��裷��<�>�1%�jz���p�s�V��H�h'����|���`��	Ί���<�E���/Lñ�4$-�8z��Z�Ћ^H&@���}�؟��B�+�W녁�
�f��L���ٶהSxދ�'C$@��R�7db%u�h�uwL ����Kp���("�j;�Q��|���u�R�bdt �j\s+���e|�[�j/s�}@��.�)�h��Lp��6nO��1é$9c%;8R;8��}Н�D��*��(Q�>K$���׎N B���L��.�������e�\�E��Y�E�{6|��Q��9w�,�TJ��Z�4	2 ��@�%�"hn������M>�ND�%��ٷ*�ֿ*&���k�5㯒�\�B
}�+7=����&T%�2�Z�%��#�_�l�驛cOW]�b�̘<Hf^�Tvw��>�S �R��ytS�@T'?�m�|��d56�ݘ�ퟩ��%�P����n�{�(�l?�,�7x2Q�*��Q2A��Vp��R���W�t~N2b�M�'�d	�M(����8���D%Fmp�;�c�S��i��\(����q7c�ֈ���@;�50MQ�7��k��Ho|.DY���&E�2H�l����;����i'�Ǝͷ��-�����鱀��ï����\9q:a�O��,Y����y�h����|�:�ml��[=�j�P���s���ڷ�k�6� U���2���29�Դ,����o�h	�]�6H<�����叙�Q�N:���>P�x�����wԃ�	"����i���i/���d��&��?�,��,�w��������M���@�{���ASV*0����� ��Ӗ�+�A��b� A�%�1�<��D~4��Z��U�/|Y��K6��P��B�r��S&}�L�"Q�KI�c�u/��-�v��ګ��bB!� �.%���s"�0E���L��C_/	�C����6Q����n�F%������Ƣ�Pt08|*I�-��WA�nV�]v_��D!=�)��x��jB�˿f�ܟ8[a�#ۉ�m�K��}�`���a��#B��i)G,���)��'�rMG����ccȸuL��N��X��R����#����,�4��n�USr� $ұ˿�e�"t�0Q{SNE�#�;�h,�m ʯ)_o'�X?�t�TfH�����Ћ9.;���a���Fr�@�}ݑz7��Ơ��Z��P�N����_�V"�E����$��Ð4i!`yPHޤ���4!蓡,��`X?���~ނ��տ�}��GL
\ �3�Ei������`���I3��sָ�܌�|I|�G�t�{]���i�|���%��&#���<ĔGM�y�wmK/}��jl��p	�UŹ7�V��4�4�9�#-7�����ゴ�X�A=�3��;��o_�G!�t��̩�Y����w���S�A�PnY��6<���~ �?Sfo!}$]����IL�@M9v���;�A`ݻ�R�'�����3Y�QJ&��gN9��KRIXŭVx�#t�ܘ����*mf�)�ϐ���d���U�֠"�	ؗ�y ��i@��2��F��}��q�Y*T�Н�rٵ�"�tD'�T]@⎙�U�ٳ��yJ	�H&���K	�҇=,��2@�|��vx.Y�=�R5V�|q�~��{y�8��nE�ɓ��L^5�p���r�?�i����naX?hu�-�Я�._�)��MF���.����@���c��������o���?WAʅ�e��C����Sv,�31h>��-ROIC����|��1��A-�;��՝����$U��r��J+�*�6!���#��>�M���U�;e�m9'1�,��h�-4�<��L�(8;T�`�2��'5T�^6�T nب\��6�)J+�#����G�	5jS��^��B9=���Ԛف��� THͧQ	+ѽ�k��������*�Y��r&:��"X����JôY��D\��8��Ղy�$�`ݕ��,����p��	����q䉻h	�G��c�*Έ�V��	!�->�х�m�]Ǻ���J�h����jX������k�\��ڟ� �)L�&;#�W�{D0TE�6��;vOt-�`�J5�}^�f�!�&!Kul9�xœ�5?�1-(|7����'Ŷh��6�;/��{BL7`o�Sm҅�e���p����w[ğĞ.Z��4�e\ ɠ�E� �O�Lx��z���~v��VP-%w�i�I�/4HC��K�:��U��x��"���������ʴA#|%aP��Ö+���3k"�z���������s~B�$E#J-$뢝&����ː���6s�#��z�cE3n�K�?���y�'0�xY�#�������o�v����Zw+����^�g!D�)�n��(����Yk!��c� ��1�	$w�Sg�cNV���(��y?�:8G�	^Uw@��E��d�R�y���k{%0E���,���N~H�D�6,��U�g6e�*�@�������Ϋ�ę5۷�]��S2t'�-�V��n͓u�&O&(*�������G3�c����V/��3j�".��j�L�|e��������,}^�u� �H�$LTk�ׅ�M 4�P-Z+��9�y��^g�Y&䮻;�����F��F�c[�^gn�<��� (Ќ��WiX��@�qjz��m�&�Lh��_,*�[� ��$�[놞DR�G�s����:�=$���7n���[��۩��Q�޼��BsC�Şc�ּZh)����{ܯxG�i��i,ǹB�N�TW#ؕ]�X�o����j���/�E�ӳ���
�/r��`�S*	5��~ͅc�4T:!>b����+��U���!c�qz��� ���l�;S�@�
�t�©>��}l.Ka~�'d�)�{ݛ���Ņ#��8O�'��<F��!ǩp_s�l�Eg�Sh]����c��n~�Dk���1��]�Dj=��S�f��<�f��?��[�b���|����6�Z�D�>�ؽ�AZ=MT��E�m��K=42zġ=�}��@��.qG��!���￧Ho;�uq����eTp�������]%Fs_
�z�]�zZ�w��U��q�������'=��%�
�M2�;�T�GGA�p�ĺYFJ�/56��9�k��M%AJYm��"xr��됛Pۧ��i��lKv�>�FD��mzP��	;�c�|�i�H7}`���O(`i�(�<:�-Y�y������,��Q����R�3m�8�y+�`p��=��N�"��}�8���dG#��o�8ܛ㗆`�]&�+S�\;�)Qof�U�0���u=|:�]5��]�vMgi%J��X�6Fo{�A�A�"����~��~謎"Ќ�2�:�ڂ�w /�كǬr)'F���ħ����� L&��U���M��::f��k���NM	J�.�U�J��ǡꄊ�).���n�F�}�"�}_0��j�E�Mwf�Axʗ�דUؖ�S�|�&��,t�қC?�!(;UQᶼRt��Ϡ�I�������#����o�J��F��Pհ��/�o~/��R���#�ϷsK����y�ő��F�g5_�Ɠ��{����\($)T�'�?��\�(1��M.q���GduB8���t�>��~g�F����n���Găl����;
��S��{�ߝ�]{W'��s��թcu��ڦ#��.��'�p���*R5�v�ml,|^��`��l��q�����×n_�1*����p�J���K��0���i�4�"^65+X��1A/m��=8���Wj�h��q�R�ShIji�}!�9���qnz���$�W�����ySc���/|
�#�0>�>�������n�
U�-�Qh;=uD�GH9A���fjF�Ʈ�Qw��Y�fU+�P�S%�-�ay�D�d�ܧ�����d:�0<�j�4����Ԗ<9z<��z����he��~3��Rm��-����yqq@���CU�Xs������lʆP��p2@��k�6���L��2*P��锅�@�x�x3�q|������|���;��s���_����>chj�}2pX ŋ� ��'8Z4�w^�����r�z��CAd��"9ָ���0�U���xx��	"'{�� 6��X&l6ſ5Ɂ���a/�Ϝ�q�+�+�q�^d6>j� ΂Y�pU�2�~IY�;�2���Dq��:�}3;l.��<�����-��K{�U'������U3�{�Wu7*��fB�W�apִ�L���=�?k$����vG�i��c��՚*�����:�
��cn�N�X��׊+w��.err���,`l�wZ:z�l
f�S
YI�����F _�KV�l�x�4��$���b����h��;rV�?��(��T�(u�7�<���oZ����s��?:<���G��}9~+�"#�Vs�m ���!��φe��;e�b�
T���+#��S�
���ٰ�pS�0+G<\Md!��_��}�*1����E5�}���-�s}M=��:�d�Fv��d��B�YM�g������щ4�S�������Ybr_@!Q�ƶ�=��c�U�����z��v��a�U	�M�h�$41d��WXE�*2�@c�(>�ONʝM����F-x!X��nz:�ʸ`�}��2 ��>14�`4���S@ۘC���Im��`8#��y6�p	�n�I�WV�/-N��-if������(�i���Ϙ���@�'��	�m�N��m�� �Wgr ==|�ȿ3�-6t�ëQ�Oۘ'�0S��}�7}	�oC������i$k=�F���شZ�鐜�d�T� ݾ���N��=x9�P9<yg�x�Yi�������Ə�S܀�q/����l�Y�-NL�q^����(3|��f�Ք������R��Z���Vāq\�N�Vj�!>�xS�*�0�
5Z�:yL�Ȗ[;�e������0J ��˟S:>^�q� ��/C��W��u��{<�]9��_�ʜ��pr�I���#r3��=�v���!�`��$����D���E��2�8c��G�R�E���kq�U3���m��9�%�����׬� 8�4�ҿhL�R��/̝>PSH��ญ��*�v|f��FOl˦�{�8$�b���-8�JE�Dc�T����a�b��@ȕ</�YBJd���~�^0��6Y\c"O�b��gIA��!�*����q�j�s�YJ���kǄYk-���4��R��ʉ��l�5h4L=�#�Ʒ�ڡ��q?lQ<���. ���	x�
�IҢt�Ŏ9���aj' 5B����L���-��$� �w���~Y3;����."8燗�s�lM[\���8��eK�����B�4�[�4�]�b'�$3�b��9�1:#�u����'���?�fo0U���\�uP3/`1i�m���N�Oxذ'*h�r�˩�F��z+e�$r�Ǚ����n�#��GU�L�2�`
��yleH)��;Nn�	&4�PIKus�&�Eքs>~�������;�`��)o��/-�wUsy�+��R�t�k=M�?�*��5pOb�<�vAFW�$�`�5 �0����g����ݓk����� �e�p�Y����K�Ð]����j��\�>�h/��w��ӨWwP��Z����Ǳ`��+WDS�"��Is J `7�ZW��9w_}��J�����R /�g��?r"t$�U����;l*a,�Nr�*�k��!=g��R0�B�X刭墕k�D}h#�!���������0����65���2�vjMu��q�:��ΠB���|I����|)�i]�:	�����}����Ssyn{��D*��%ZL�й�1؏?��W�1������?���'I�ao���#`�Q^�1���W�_�A��2�nc�1;H�kT�;RNv�p�|�����ȔY�bu$'j܃Η��qO*(��8q�Rp�lK@��M7!'��C���&�yp���\[�y�.��Zݤ�<э�����K0�H^�p A�x�G���i��$$a����_]�5F��9�;"a(����ۑ��bBti
�xU�zC����F,�!/�2k�����
�4޽1s
U�WJ���]��t,[�����Ρ-���i�xs�mWR����.�]/���*+�3��Q�)9�}N�]� ZhR��������My&��
!<�s�
��>%���+����4,�,�@I�W�&�$��4K1��r�h<�h3:k�q��iPĥK���t[	�_#,���f
�(��hU��W��ĺ.B�@ۍcUTف��Zд��������8��K�����&��0BIY>�c�;���ME@33[OD��z��r�3��ބ��"$�w_��yu�9q�#���O���������h��ٚ�C�L��W�8o���h&F�����x-���es3�D|H�H�7{O�`'��
�����{�uY�+��Go�Myԥ��+�Ru�r�,��>��f�@MB�/�Yx�j��x�pV$�
9�;���K!#�!6̫�{'�<��(%B �%�<�Z��t����}g���0?S�a�1{�ô����5Z3�P�.�>m}�q��ۋ�-ݍ4�iF����fe*�X
I^�u�_$Z��[YѮ��P+Iv��r9���ۺ�$אb2/'+���Sd)0�͵GK�\i/8���doT�rj�!'�Gɣ�isBW���'�p��ȩ1WM^Cu�'�sfNl�~�+�A������=ȫT̻`!���Rd�m�����Ƌ{�!��|��`{��J�h��c��`Ij��~'��m�!��4�c�3KQ�_� ��j���}�?.��n�,]�~����]Wu�-�,��N��\m4��+���s�(���W;�ğQ�5�P�)'��:Iq���eF^��:�])��Y�vt�S��h�,?]ô؈�v������z:$E���I )y�ƍ��3e0)�R� ���0la�����r��Z�{r�����4��+�`���z�A,���ϛU�Aa����Э����тn(�E�̧�71�@-�NĆ9�&�;������Dѿ�>��D�h�C3O�O_�$G�:�t���dO7�z��8�i��m2��Y�Q�b0x�r�U0�  ��������T4�nS%� HX2A�����>Py�8��r�W~(}~ᦤ"Ԑ���M�*kGM��%J�9ڜ7���AHB�Z�9c�'l�%�W �(��*:�7CT�,����!K�5 1q��W����H�b'�r�/�vc}��9����q��n����0��jёY����:�k�6;�
'�<t��� f���N�� ���i�JO�&�!Wm\qE�hi�{��˰o� ���-�a
Z���)�����@��p���ze���8ϙ���ϩ0�M��A����%a�^�o��A�[�"�9��S���/G���/��1�c�ھ>o�;�v����j~�Hf ���D�*�_�~�Xpxl��T{�,$�����-�¹)k���7�x���M�M�r��/ܛ�uc�RɎt��m:FE�~�Ջ��0�j�|��ֿ��}����zX�-��W��$F�_R��I��6�d��z]mE]��V���0:���U��\��a���g(�S�\��R��sGz=ڭ6'g�O�F�+�3�it�`DW�Y������-%3�̟f\q�G<�I�l�����(Y(^���2�R�5�� �)�͂�NA�*�H�7�7���E�U��Z>��4�8�C�0�_�^㘗���Y����|�=�i���ء���(l�ҽ�>L���?��]�l)0��Sa��<6�0{fEP���� !�p�)���F�;��i|�F�C���vܟJt15�BQ�ϗT�������
R�?lk2����@o1�%�a2!��(s�@�:b�o��F]ñ��8 �tGDQ�<zK�u�*M@G��@7�G�Eq�y�#[0�J+��c�l��="5Ӫ��7���K9"%���n���Fr�Z�1u��q^�
�ĺ������*����m Ww�@Z�<��t%�����Qe��9���vI4~r�@�:Ǣo�/&l`�dɄ: uA)��7��Z��}�Nxdݼ~�֖�P@ퟠY�u.�*��������bG9�QQ�,�AN��6�җ �j������E.��m���E��p���y��ZDv�#U�2|D�������6B.���dүحQ'"[�M�к��}	l��X
�E�z� �ͫ�ʮ�KV���P�՝�k=]�/Y���Ջ�3�l����]:D��)Kݠ��tC;AA@H���L�r}��
n6cT:���*+��F���'-�M	;��Ų�����L���P�l\uD
��oo�F�v�������͸�G�M��s��q��K}�~�.//$	���q���m�Y�����Կ��@@ɹ?�%�n'pչU�"���G����?J}2Ja����}��/�����5�}�u`��B_��)��H��)���B��m!�f�D����Ҙ�jF��Y���W���T�_��EדSq�B�� �e9A/�������T]z�b��%Y]�D�������9�;��i^��چ	F7�x�͆+;�h/<���p�zõ�:�G�~('?�s	M�}����s)7�������Ocpf�}�<���7����dɗHK�$\�!;�ܦ�� K�䆏�As�4�L�TR4J�t̕����������"�H>W;I+w_1k�����w8�4g�4m}=���Y-oI4�lq�f�v��%�9��$9����Ld�wφe��Q�nB��'��)2^�5R5��Qa�k�>ve���*��ݝE[�F�%$�YŜX
5��Ł�����QU���v4�;X�Wj��i�F����H_?3�Ś��F�~�s[=�&yR��|v�5a-��*ls�
���=���&37o���Q0��������i�dA�W@�����r����J�Ӈ�I����!ՌZ��VTDZ��o��b�V�OȐ���r:��>��wp���B�4�
�\���Ȅ�Y�jMkgFs��[*�1��ՠU̞i��Pl�P�?P��D͛�Q��,��JQ��K�oY�+'nK����D��Nd��Ř�+V��6�<һS��;�J����*p����*�4���5�σ�� ����P�������+�v����5C;��F���;���K�c�.�g�+_�^�I٨�bz5A�6v�'/��מ|8$����� ���ped�͓S�W�j�8�s��=�2��&d5��-�2�r��	>6�������.�{e������CfC�3���ͩ}��W�#Ȼ�G�R[����F�y�g �tj��6�^b��QW^AY��y�51�HSP��΂�)�L��Ht[���4��͚� �»�Y��[�s�"�������7w�����PL]���߇��-�ӄm��+��38	�3���:�W�},�x	���ݾ�)����6^<�rr{SM�H�E�>>48��;��#�h#�>�pH^���F@[������y\��+ ���$�#��q��D�>k0M�;d\�y�[j`�K����}�'�N)l�2p�Z�������"�";})�z{+��:�*%d�Y���V�6=�A��/\�7��9��� ԝ}H�����Д7\��?���d���L}LIϤ=.L��<��9�w�Պ5MuAG["�8����;��kw=��*�8k�#*��T�h`d�����*M���˫���O���2ˀc<�e�9�ÎP�H�Ø�h��w,e?���?_5�z�W�Ύp9aΩa[�"��{�EE'J�E	O`ᝳ�S3[�Xޙ@E�)$����2u���7*Nƺ?j�W|� ث����3���@)��( E�-Wqe`�C����l� ֿ��d0-RVk	2��ͭK6�z�X��5q(�4�,QXď�=9�|e>���\��f�~�v�-rM1�������5�#VD��o�ګ��@��UR�]{I�,����:�C�'V�R�h���o�M0���n�?p� mD����[�V�u���!�H��?�:�\�Q��Ohʻ�z�D�c��ʎc���sh�
�|Iٮ��z��_��O��gt�5����s�uS��I��y��
���]<>���L�.����H��j���Ί���"� �=?�j��sSA�}�Bl߻���q��/:��9';�OF׫@]�sM��=[���@�=���_�LC�������m2�,l�k���_��iӫ��wZ��w^�@�S�S�¨hf��7��)v���6>!DS��|�E�[�g��Ba��+��W�EL�6YP�1�ml���Ajj����RD7����haZYD9��J15R��Bag����ݖ����Xi��T,�|{�:��AK;�^f5�܈�1�X,�j�х��| 4VWDP�faϨ�k���"P&����x9��n��C���Z��]��䜿�o���9�P=�1����RǛz�pb`��Y~���M�06��K�����ˢ�Y#���	�[9�
�zn%E�J���J3d����[
�ix?0R��VIBP��U�[Ys��EA)a���!MuՒ�|׃@9�燙����4xl�844JA'Fy5�o]O��$���=j��,��A�����&-W�$�S�ҭ��'��_�C��mP�X��K��8c���`[�U�mo�^�2Z_�#��6�k鉱iwt���'� =�Yhq=$���O���gM�Q	����F��m��i�>�w��5^��
rV�=%�)����TA(��ez�?�*Eɐ:��2���/>j�0����֦u[�>�r�~��ƭb�n��5ݎS�L-����9޾XF◂p���_��XE�A0�#�����:�b��nf˜�����|[��YY�=O���/��Q0�ϥ��EfC{�d��)n�T6HO��t���J@�Ȕ	^����a�K�j-��	l���:�j���u�C����%���=fqV�߫���_�{.�{h8}8�Gu���d@�G4�w�<�ռU��~j�LM�=֙c�fS���.�O#;����c�X�]p !7�-��P�Y9�@E{�V�EuA���gi#�6j�C0�^�ے^�J�+�8��w���e2�����Ԥn����*�y�Lp U����&AR&�,>�|^�}���gSih��^�+��sB�j�+��[�C2��Ǆ�S'>@��k�F-�[�W�wq_b�j��y��M��a��	��c�U�����{a���!0E^'�`��ޒaw[K��(z,�s��q� �t���\s�;L����Y�!���d�VN�i-������:���� ޅn~ݲL���ᄵ��&�Q���@���%�ǵ�}�yEJ�)��4�(����HO���=ݲ�r5g��Ș�_B%@o���K_C��tl
�<e)ϙO0����1��?�E�hM�9x	@<��aW�l��!�qm��_<������!s��q�Ll�ߣ�D��uG�S[���?�V�e�A�#���C�U��z���.O��	G������F_JT��4|2��N
�P�br�
e�z�=3�W�.(Q�pC������Kz���z���ئ�d�E}b�~	PrA��f������v�W�����:y|͡���ș���:�nU���i��\K����Gj+Ʊ�/����ҡ��4�Z�稔W9��B�'l��=�~txABCW�8�pc��;KIn�+sK�}�6Wt"q�E�k߲��g��L�`�-��2���q٩��\V�G-� 1雂͓�������<,�5������j��3N�k�[KE��s����񓠮�ɵ��M*�ϱ��������R�]p�,XD�ҩ�R���2⦹�ɴ�W]&KI�Ƞ";d���?�C�mUi���_]� ���U[��w�a�Y����_*(�)�������%�L�kF�%fS��QD�w#Q�d���𱌉����yS�Ө1kV ��s}��e[����U���C����=XX�ӆ��T
�[���O�N��Mh���/&Nդ��獫q/x�o� R s���i2� B�I�DK�i��Y�4�tf+ڕC��!�L	����.$��X/�kԟl�����q�!hq+ı�j����K���kZAw�*��
NPxe��GZ�3�EH:��
i�L=���#���/��R�~J.���Ϟ���%&���֎�����w�%H�A&6����B�仾_A�|�\�W���!j~�"F<�"c/yd��-����J47cu��ܾ;>aZ�P*)�y�\}�^�ʳ�N�Z�3pP����2���#m:�p	�:�����bFX��#�n.���?�}�ڝ�����R/�����@����ӸG�͉sp[�S{.ӱE�Wѭ��E���'XԦv@q3_T����<��w%�WwfX5�8�ŕbe�M�Q���b�k��h�8Rwi5~�+g��=H�� 	S��@�F�����P��x6C�6 ���Ũ�Rvf]��h�REo�sPb�r�(}(�� d��?��](Ҝ�X����r�~z�|^k���W��{xo�
��V�?h9e1�4�eH�{� /е��s�VV��� �:�4�1�ɚ��N�/�v.	r�O��a����_j@�o�0�YK���5eWdMb�?�,CJFo�g- �a����L2�jW|5�ZD�kB{5u;OT�<
)Tv���K���:XHܓµ)��N�e�.���qS4#�'�x����y��N`.*�s�b���N�����O�6r!*0+گ�p<�'�恑7CS���jӽ� �E��lX��"�a���()�TQ���a�A<�|LÖ��Aj6H��{�.�q��������4�h�|�1���Ц%�,���Ȫ���Bӟ��T��9�USz�y�a
p�����X%��I��P9�H����.�]��_K7�)�nݓz�9�_�+�7][�ycvȎ�����`H���_�%<�g�쩃�6/oK5
�8���_o����i$<3".4Щ禁��r��������6!�>�ki+	'&B`Xn��+~�n�J!�����c���ǮU�����4^T�7�N��m���'��|��k�!NU�3@��&v<��È Բvn�s� C����?�e�ʄ|��Ҽ�[���&Vm�[��/M���}��0�������w�{��Ci�=�1�A�z�����3�0]�t��_;o���N�0B��~�xBWOTw�����珦�����B�&��KQ�Z>�Ii�4[�C{�V�W^�`�&dA�vW�f	��TF�0�2`�����(�l��LNi����n���\iPKkE���|��c,�x�(:��=���

�)��E��@��80�b�Vw��U:E4��V/�/���z�<t���Ҧ\�ɥEŌ?m������Nf�m�Ue:�5�M��Xq�^��]�/\+�Cwֳ�>%��gC̡v��(y;���~���knr�q����'�]�ŗB�ϸ�t�S����j�������Ҵ~}{��e���(��/��V [I��3�� vE��j���v���h��+nO��]ך9 � ���|�����肕y�PI���H�-@��I�*yC����U��RO.q"ӯ�:��w�����W���7�ë4Ďt���K2j��A9}u�}�$QɅ�@Zs
.�85�\��̽���$�Ֆ��F��I�{ږsC'������(�\��#�� �8��*H������R�y�^*]&�F(ZB�W�_D�~iJ&��bփ_׫�4w�^�xiYbɞ�o����|��0S,-�,�^��V�'CYP^U�g9��ɣHC�(�`'�[�#΍��K&VrS��y����ϳ ��H�Ӹ���m��~��S�{�䓗��Z�s((�l�����XZ��8��ez�̀�I��.l�oq���$�P���sN[���]�@H5J0��fQ!.Q*�V ��5�#}/X&�rI�פ�)������L���N餝E�����m>�����W����
U�A��^�������:A֗����w��m)u%� �Aڥ�o���2�� n'�:2hs�P����4�#��w��*�:��p
�_'_�{ɣ"y$��)���I��{�M���TY��=�˱,V\�o�w�m	`9B�9,�����|�F�;�ן�X���Ύ�j�8
C��ؙ�?pB^��k�;�G��7��s��#�Z(����۷���G!���{�f_��|U,��`z�X�|�ۥ=+l�4t?�흈F��'�~�ԣ��\���U	%�q����с�5�YG�]H�U�T@ ��q)��~3��L���F��t&�i��ϒ��!%�LbrV���!��s���c5�n~�;�/F�Qo�pn��c���'�L5�3h���0�R��{�%���Z�ʜG�����Y�!x#����>)F������E�kPm!�C���R����0Y�~:�=�E��";�7�M���.@��;���aVw3w��G�(Tb����$���Đ�$��m���f�%��P��I� q{��V�7����!V�d{�� ����m�퓳������f����ݣ��)�fޜ�I5�l�
�	�.Aa�I�W�v5�wHUO��~vP-%�cl�*�d�u��dn��~�_���:�����.�1+-�pF��E���@:��q���ur�ȟ$������n����?$�+@�d�vB�W���᝱ԩ���?�Dm_�e���g^��G��p�Y���:Uk<�7��w'��%k� 
��Y�?�l���h^�kq���	Ocu8|�I8�}`��U|����řd���f6�!m���_j�˄�/���6�jTʏ:u�݇'&� v����$�@�TN� &�	s^����
���ihve{2�~�D]	��zk(Q�⿁`)4�J-�c��Y&x�JD[���8#�|�8�E��Y�*��s��ѭ|�ؿp/�k Ұ\�3]�)�jʈ$F���$���)NAI�e��;4��1<�J���%�[-S<2NN�)��=���<A�|����ru=�>�֠F-
��g��+���6����!�g.XX�P?V��nY�Se�~�UG=Um��bQ��0l�����֬�*�f[�K��Aϫ´M0�ݶZ��dQ2	��oL����'���Hy���R��v�v9y�D��!��e�P܆����Vxck�E�Z�N��Y� 3@�4�!Ҧc)Jő��޾��Ƚ�Q(�n��/��H]�>���nq�J��|��M7�վ"sG(:��<V���3�o.g�����t�v�8�Æ����ӥ{j�wd�yv���K�@�{x�"D� ��|OU��Rt�0%�\�r��M
Fco�x��f�3Os��șs�6������Cf��>���N�mG�}��S���qD���y�6Rg�h_�����d�i{����S=����'�D�_9\5 ��Ԅ�X�{� B����ռ�Ѯ)��0�ǡ<I~_s� �* ��c�[��=� �_������F9Fߧ�ǻ�
J�|Vd����N�J�,\�P� ���o��R�@�WcI�W��� ��F��H�Ű�{?��b�q�"۩�J���1Kރ:�B>�1�	�G�+���M�S|��k�K��c;!����J{�h�n;�C]yl<����Y�n]���b����ß�2!�����Ef� s�gB�Pg�G�-
�Gy�Z�������c�Sa�U�K�83�⳯�k��PuAH�T6X�D�L��KA�r���#w��,Kc���O����֍A��;��o���uyQ�c�	;�Q�lx�fz<:~Kh2����>t����|mGǓ�Ą�#���y�!-��K�҈e��������%m4675�s�)��XjS�H���GT[Ix��:-i���zοECP{Ԃ�z�'8c0M�
[~)�
A�h:Lˏ����S�(�gB*FW�X��@~isKg_����zY���' �B��)4C!�) oW�9z��Q���|�2�]:3$����B?�,�:L������j@�&/r+�A9e�ﲊ�[3����p|����⓲Ό�g"�$�Ѱ��;��?��Z����N���@Eb�@��uS�]�3�~)��f�C�(;��x��P�!���	/&?���sx��Z�4Qԩ&��32��8�%��1c'���M>Mb ��	p��`�N~+�O���j:�w�N�%]-��U�1��R[�+S����������X�|�ǡ#����-iH6E�z%<��[��9p������ I1ޞ�-q�ƶ��9!+���;r�}k��Q�n����g< aW�	#̰���Z��w�+WgYC��bd��z�ҧ3j���_,�Q*�@?.ey`S�FWqT��$�(�P�ȜX�d�NDk�?K��f�X|�>��?�?�^�148
s�M`���Ԓ5���8�a��HD����������4���������&~�(/�B�~e�0�.�Ѣو9q�-V)9[A3,1@5�ʋ���>�V�H�s�r �w�2Ɯ�/κ�i������]p��<��4ѩ�N��������))|� RE�P:F����Ӂ���d���X����%h��#f��؎}5��bD�h�iȌua���M��,����Xc���<�U/܋��N�aV+�r�GM������@A�Ky��oP�d�vn1�.��8'
g,�kͺ����hE�D�:��"rHȓK����M19���ZrQ����ܠ3�����b�Y"K0�v�E���'�~Z���6�=QrDVM5�fYB�Z��H�X�Nڌ��d[�����]�Q@$pc�Q�;���x(â2�f�ׅ�����j$鑝�r]�WE&�,7������q���6,�Ƌu+�^"��%�	�g#�;��>L�/�X��ޡYAas[z�2[��v�����YB�t�� "��5�Ȑ��vFG_(	���"<��SU�d���7_����k󄡓k���Z]JB=�^/�����o��a����v�(��sU��pU.���[)��F�C��k�|c�M��#���
,�������	�R�%o�m/� .��ٸP5ͩ�G��^�v�ߦCA��7�]d�x8>]���P8ú��ˉ=J�i���OM�FEh ��Ys��~G�h�_Tx�M��|j�Ѵ�E�Fxd��i}-��y�'\g��J�f��v�z4�g���TD;��%�˱��!aWѣ� ���a�F���߳|����~�_Sau�q�<���MZ�h�"�&a�(HWF��[��4B'�x�8�o��D�l_~Gy$��"H�����ˢ �r��0��:n�r�ްmz�W�y�L��l��5Pσ�)�%��v�6Jљ�z���)�^����jھ`F�*�Ͱ&��xx�u��v^�?�?�K���w���V'請U{^m:tC�o(X�����oM�H�!�m6�b�ۀ�n�"ۀ�{��^A��t��T"�r|��p(�k��Y��~�lu�cV�X �З����/�7�k���\��/�/\ĞX�7G�M'rV��s��[���$�K}���Qv<��Ջ���Z���������@�xNQ_�-?Y�k�/B��[�9��/����j���X��"o�_�w�ڜ�6��5�΍
Xe��̍�,�e�n�Y ������+i���/6��Iv��'�/��	�h����D"z}6ɡcP9��'D��_�;��F�Q`��Bv5��}z9�,s��Ju)`߃�Dy���\r��(p%�U�<��Ѣ������$T-!���+����%�[�;I���+j�'�ܝF]���(8��I��?��5��=����j�N�k���A�R�H9)l@�#�{���ϱ|�V�刯�C�(}w�|}��ϻ����N'(����bS1w�,��87%#���$}�:��cn��dɕ��"f�L�Z\h�{��%8}ow kM��eg��Y��Ƒ���H/�V+�����)��o��v �j��c4���zHq�Ϣ��g<�o��x�Ok���j���Y��l58p�ޖ�.���b����O�C��@����	@3q.�|5�qך/�0�!���M�f�	�#�'y՝���\��l=�h��0P>㡵�V�{�{Ǽ���&FS���/-�P�v�V�xF�w9�/��A&���e�U5�}�c�oY6�~*��Q�>��X���)�C���X��l_������иgܪݵ�]<��7�
�Z����׏���^�G����ᬛu��v2�3JOd"[��(N����Ja�=��Í�[N<m�L7�(ii�P?�#q/p�69&1�#9�E��r�R�J�*$T� D�i�8�6�ZYX�!��ϒ�L�p��{9���`ɏ�z�\Y�t��u��]ҽ�`��vF�}��ᔸw��L�d	zr̰��a�i��b�)T0����c���{�n<�&���=��:�=����`b�:�#�k����bAG,���=�[��j�	��jS��9<�3o��L+�R�
�ĵ���U��"��-Q@a@�|��f+`7��ս?\R>8}($�`e��ߙ�nD��4�O�lyk��9�Ո��wT���s�0��v�X�b�NP��Ď�47C2���[!�RW� j�f���Q3W@���>�WU� �6b�"tS�M�i��E�,��j}#�<���������SK���1�s{��˥�6M�����8M�RN��P�Y�c�)ޢw�ϰ++=����/X���6�}�T&�^Ӏ��������>�<��x��F�T1$�E�����������n��aY:��WV��y������.zX[r!�����{�{8�`�bN��(,�x� ?`wfY�̦�ve�)��-�~]\j۷�
~�o���l p�=g�咷aK������v �LMH�)��N���FM(μ�eN��o�w�+��_��Kgp�.��Ue�Z�pץ1U^��j�#�����8�({I�?��"T&�P~�7jZ�۸/�B�Q��r�K�C�	�D�3��`��<d�rD	{?%`q�4V�W�����T���X�����3�n>#֩����J�����]�L�b��>�l��3���HR��4��1T�B���y��O8ΘE	��l|�쥎�$P�)'����c&���̌n�G�{v[�<;�����
p�o���~��l 3���j0��i��h!��/ ,�P�~��NJ�L��o;8���J)� j1�]��}9�(��"@.`�����S�,����4�IcTC`�B��15mP��>!xF]	��q�������S,�Q\�^���u�����X@̋�*�A��<bY�M��".)�W|�����U��/[��R�W&Fx7���;'�vi<��Jq��cY;>ĩ/zy�q�� ����D�A��Nu�D�k�X�X'���-|�Yp]��ݜ��rt���k��J�U���*c��=�l����S�h_dq.��qj����"3��:�7J`����8dc���|�7y>@�ན:�l�y��clg�*k�m�U@������G�q:�3?ڼ�:�C�����E�"�X0�RS�隆�@e*���y[`N9}��E ��:}�h`��*f6�I���k���\��K���@�_o�����$���o����S��Vx\d2��j����aSz��8L멵c�Խ{�8��µ�f�j��r���� ���+����E<����;�s�r�99�ܑE���v��>3����6,R��s����ӕ��y@]|�{)��iy�0J7NJ�mw<0r����|\qz����*�Ƿ��;¼U7Ӑ�Xޤ][�|B��!@�����Ρ`Ij'���g�C�s����'�4gu����\��S�u�=��k�9ػ�-�a��U����U5���'�MG���k�̱�ԋ0{8���ԝ��Ű��Lȳcb�X�������"�٨Ʒ�*ᫌp�b�'I���$"�3�;�E"���F>��,rni�c"I���qFiL����:,�v��L.>�̂��(��'��r@��Hv����I��r��܈�SkX�mS��x*�~[��:�h���]z�3]4���V���3��o+���L��d��-�*n��`��x��w�����_�VV����x�_$�i������2��j�a����6*�B����;����,y��t.Ԧ :��'��f;{��˦�e*���z��vO:`a���h7þ�����_��#Uor�5���L+�&���g4)9ɐ�#~�=ܵ��vl�C���aGlk{0[^�y���"���!�2�C�|`����Q-@D��z��l�L
ƭ%ʺK��X���ZX��T%>��쟢��]d���!��q�UR~�ݎI�"<�X��P@Z$�����+��1�j���h�L��J�\E��v@R�:�f�v�}���=�G�g7��������=u# ��8n����[�QU��+&W�-�T��9���;�EAY����b����)��=�L�z�F�ԉ��P(R0S׭ӹ��v��'�`G*�\v%�џ�;h3Lۄ���?������}�I� ���󥍥5U1>v��X{�,�� U�c�kaP}�R�aC�G���e�bg�^�h�*�uAGPb��z�H���V�v��)n��"Ztk��J%r��N��rȍ%,o9ƀc�1e��,�bC4�l�������;$oyL�qqR�v~��v�#�Tո����e�W�_�`R޸^b��	u�M<�Å|��l����cg����@%7EHaw�B�vF���3�wV��[w�cs�/^�畒��~H{���%'.4}�*kBI�G�9��(z�<�:�����r:�#�
�Nq`�gV`2??����*�=:�^G�Uܫ���iy�DVG�e�V~Sn�daXk�mk��Ų���?�K.+QU%>�<[��rL�a�����0���Q&�z4-e&�-�j:)D�}]tǃ�Uk)�m���R�p�!��JN;�^	.�uWX6�Sj��P�B�Z�\��ArtY5 `�̑U�����6~\Ep4_+��C�K1��PJ���ӼD���J�W���7
|T�=�&\�@x��V��\������]���S:E�L*(긁�@j4��m����QA�ܪ�h�p�7Ē�����QQ�w~����QH<������^̿��2�8��__ô�����U:��1�PIP��h����f� ��ګ]�J'���qy�t|�e����4HK�����q.���������܎atka�Թ��G�GrN��y]���
�|1���UM�|��m)�]~=���0xh�t��:�4m^I��h&��y�<�?p��B\�g��e�E���r6��+/\Lc�D���|��3RCaLf�52j���@U�������͵�jϮ\J�ٺ��W��+���n��V��,����1���^�i�����{<	~	�C�]��k�N&�//#m��v!l!E���R���C��4fsdb�8��cj���)"���n�"W�i�/�S%s���c��/Y݃���j�Y�Q����*��/��=��&�|�'N~�8=��{�ԄRQ�̚ \��i����[e�Kg��v����±��qǭ>m^0ZG���p^�v��v��4Uߚ@�Hq �����{?j�k�9E�w�M��jN�D�5�v�n�2
�?`���&NZ�Y�js
�E�A�/KY��>�c)A]����ѳ���U�X��Xu�@��Wd�F�=(�%)}�����`vW\b��xh�y�J��$^.%�4�DQ��U�7嘠5�k��8/�*�یa^�2I�[�p_X��ؚ�#�	�@,����3c>w��C������N���+d�>T���]�x�N�L��`�r!-F��gs
Bx�7S�=ةIm�@Ӑ����� �C��=�nB�;�g8e��el]T��]_l(̼G˫bS	�3�W�@SG��ľ��T{(7iE�1q֌r`�;����B=��~�2\���8z��E��� �w�mo],~rr� B)i@܇�r_��+	m!ʚ�R�H�J���5.�l�Z��.� ��-����1�`�Ef^ ��x��ِ���|;�/X���3B\�J�[A�n�Q�;+p���-��z�`�v�i���%oI\]���F�m�z�߁����3;��.�
�z��*��A�N�Ѷf~����:K�@OE2zVk�X�,c�M�Y�b�?\�ϠĽRҺ)F/���l|�7~3/��s$d�6�Ȳ������+�S#��-!��;P�����Ӱ�G��v����Eq,yv��$e+6�ܿ�vu�	(��9mvg�ɔ@iA�$�=d�}9�����W�[g
���fa�:�!���)��{���C��/�b=�vw���p�[:��lpL�f��o:�Ȅ>bwy�Qo�a�5��1���X��L�A����S�x�cSέ
kc魱���)Cy����/@W�W���,_���h G����C4<�/(��O��L6����et0M��ս0ʗ�����,������p���k�<ˌ�����(�
K�Ջ�Sf�o��q���r6��*)$ʲ�gKzA
r�~�y�E;ɶG���v���-?�ΰ��ϒ�q9��^*$�M�����b��֍��e:�Xb���Z��h#�=�����p{fgVw�B#��s��\���a���ћ�]����U&�2��;�p�0�i��]�1]N7�8-�iP����An�,�}�n����E�1�F��PNhjT��D_|��l%�f�B���l/g��g:��,�q2$u5E���# �`}%��A�V�� S��(yH��D��h��m' f�q'A��M����Ԭyţ^��h�6J��ghh��6�=6��y��ˣ�f�����Y+k����p9�=D��D�R��
��[2hm�J�l�0B���(]d��:=���־��4,�I�w~�����0k�����£-:{ĪJ�&`#�G�Et
��:�.��4�`wv� p����փ�^{�rZ�$� a�p��^�܊D���
O誩|�<s��!�=k}b�C;�4 �~����W?&@�_$CC`��=d�%c�E=��!܏x�n��}+Az3�����5��\�#pсbY� ����8��DI��cgn�K 
��cyd�^���Ӄ-�q��I���_3��r�*�x�	ȪЄ�n����ѧ0Հn=x�_��ܼ���pMdh_�,�U1��T.m�C�oµF]�O5�[y�����ʉ~�u�xs�;�����_T}�MO�U���׈-7}�	�Q��w�ەE����B�~��ҭ1A4���u�gtro��T�!W���;Wo�F�Fj��JS:�=Z�2�u�;:
r�����RWc��c��8�K]�Dl����
=���� �?�"�d��g�m�]�r�l���V��@�Z+ޯ{��bd���𰕭���@BQ���?�U����GH;փB�<���^m%�3��@'��c:�� aB��ͦe�.+�����i�~�Ir2�h�G��?W�_Q��Yu�l��Ɂ��P��F5�	���1��ajQ��k�S]��&��*�%l���8�mǬ#�A�\[�ν�FlZ ��'z���i����8�����+�2Z����X��'7��gD�E�����ݷެ�}��j3-&���?����-�0���
?	o{��U+�� ɟ"��k �!蔲�h&N�(^��Fa!뾒=�JO�"��O]y�����Z"��db�_-��
9 ��j�x��J��!�qƺԱ&#(ߙ_Ojhon��Q_]�Pu��S�x=GL�nW��B��S�e&>J���'���i�d�����7]��cj�l/�sI��~?�6+�~$]㯮�_�+=ӗI��sf?�lf?�`{i'~0��!vMXc2Ǝ��O��:F���*��d�sAo�'�E�>[���\�1͟`,쬃A���fm�:[Î�۔�#�5�90��hU7��;h��D�s(�� ����{�甁��0��PnTv����{'��b�UH�:����&����R��B���nu�h��� ~!`��������p0����,��v�`��8U�a��?��F�����@ ��C�V�bP�W�S����-E"�cN������?���-���h��I&$�`�{f���H
��	��Սg�V�b�;��JT,@�����������ܯ ��6�87���Ş�0�r�G���B<l����]���m�`�z�������p�z*��5O~��1�@�	Q����R`<@��I��r�;���Ç������z�x�=�>�""D ��l;9���¹5�׋����x
�4���L"��꼳#�����Q%�+%hZ�~2_I���L+$�?�/��*2>�b6Ѻ��g.B�sڊ	�-�F���h90A�E~�`���Z��Գ]��㧘���:���u-�R㫩9`D{��s�����o��1�Yٳ7�m��H��m��1��_�z�Y��>��eoi���o�*e\�f���t��8�R�?<�\(3T�j���{������g^\��
���a�K�,_b��Zct�j#��!΀�RM�O�$�0��������T�����Thg�ګL}oʀ��j,�!bwY���Y����[+n]?���І3B��u0+%5�t�L lc�=��r�����G����; �Q�$��Y\d�m�����2���Y��蹨�"P�4��wGn$��3!��/y��F�a�%uh��u�ɧ0�L&�W�e �KT��z��40�E�D�8lԦ�/=OK�{�I>r�0�+;<1���&����cK(:�PS��|�� ��h���?�R��"���/��0�|��D����ٕ��6����*��;=��G��ˉ:b����A���j�x���q�,=�ͼ�lwaηe�<��",:P,`��=抖�6B_(@6G��P�����Y>I�-�OG~��^��Y���m������sM�rs�n]� �ã�k�m�0\jE�Z����[�"��#�Kx$��%D)Q�PQu�C�O��NY�ދ�,��·9�V��g������ӑXØ��G ���z��g �w]J�D�ƽ&`�_�P-�/��W7��*�I#�W�M�	�n<�ۏ�z�<�!��cȬF�Q9`"���_�l�:��l&�� J�9�._�p�8�TG��Ey�:ڽW���g"���D1S�d���4)��࢑��ri�u�����!w��?9i}��q�1	%Ntj�I*�_�$Z-��|3�}1��=��,����и�boP�S�E�
����ꇹfb�B��a'���Ô/���f}w.�Ke6Kwk��J�Q����#�_�ތT��w"�i��
p^�ݙ�?�#ܫ��M�`���o(�^9F�����{/�%� �}�q�sdQ,x��R�k;���qQ 	�R�%���M��U	�8��.�%$Ԓx��$���׊��H�ݕ��5��
H����zY�J��ω�;|�.c����J}�\t᭡ ��+���?�-���1n�v���5i�^�F�u��qO	����Ӹ��y��(��P_�Юl���7�	+9f�bs�Sc5mW�a��a?T$���ͭ��)�v�i�H���g���ߦ���>�N� �����$�B�pJ�}�KWH{ȗ�ͥ�
=��X�>#��xAg8�=:��$��[
��� �����H�(��jk�Kʷ�jG���rVJ{��g#�(�k�����Ť>�c-����5�T�m,vu�r�h�����ݧ�j<����^R[%���8VIw���n����$�(�9|�A;O�9S6$�WU�������1j���>��OL�8�ˏ.�"�c3��e����*�_��5>"���n�[��^HIA�L�ݞ~_�?�����Oq�N��$�P�X�kJ����Tzi��Y�	p+p����zea����l||.�P��6�ʥ�7�#c"8N���f6'j]ZVQ���x���
j�3q�I��'��eD%����-��D���y�����]@Ӷ{�3;�LYkp�VG�a7͞�b�ب�R�y��>�\���S˴�i�T�]7ψ3�} =�վ���y�mc�����b�Q^:M��ȝ��l������=�q#�V�]h|KWgQy��l��W��hR�:4o�r=I�ӖP?S^�*�5m��R�Zt0��-��"�y7��Iԓ��P��a��-�x�oK=�<q#�����;)���Nn
&�N�p|�O����HU�i�䪇�Ǫ�ZN���s�M��sQu�Go�RF�ob�o2ĩ�GH�73���S�g�@X��I�'��.�W�4d1�%��ۤd��C���`��h�l(�J�s���l����XaU[v��L�2+�f �=�Uw^��l4IM��/�=���C*F�'�^m�.*����+
�-n5ө^XS��x���2=���i�ev]��ɂ���W��0��g͚jð�O��^��ޚxkd�<�m���i�]�,i�Ύ^F�*�o�-o�����8DE�����Y��F�s��%�W?���`���k+�q)1~�/1����X@W�ku�b�aQ&D�4]Þ��z�Qx�j�����������^�J��16�Zm�"�UV����[�J���/��p��e��>'����~�gH$nJ��/q��G�N�'�Dˢ7�+ ����w_ײs�V��*�^��m�p�����v����]v�{~}cq�-!�t���/x�������w�]�5��~���JH�C�7s
�g��~�Ȧg����7(��Y�, ��,�����Z�B��9g�M(g�k��~C��h�7�\��ނ{w��������e��i�t�pe~H=+��Ŕ3[����FEJ�i�I�Q��B"�ꩵ�X��T�X_�_ѭ$�mˤ���f��s��=��eb+����KS�ђ�7dvc9������da�}���Z��yY�3)-7�R&���v����0]�J����<�k�[FS#d� ;����"�m �B�tDʤ{~ή�t�'�%_h��4�I�#W1�D<]V<�����aa�E��w��)���}�>%}�_m�C�w��e��	G6��̌�QN�C�Sp����ɏcپ-8� RPk�@r���t#��M�R�it����)�����v�u��c���1�4K\� ԇJ�4��ZZ]Ù�/��6t�i�!�Qoq"���������
s��A1	����{i�����wȰ�������tܺ�F��ͺ��i�yв��.�b!��z�C�6_����b-�s��l�|�m�i�H�I�m ��>�:7z��pO���2
�0<��V�Ӄ�ZW��a�iy_/5�FS��	RX�̥m�T�	�c!����Z�omQ1�Rt?p����97��)��K<蘲qi%'�z�(��l�d��%2��2��5��"�4�vSQ%3���� 9	� `�y��<}W5\옟�����C��9d`��6�슂�ѽ�@o�ms>v���B��4�1��11!��񦵐����\���w��"�t��n�d>��ٚ
�.."Qb���vq��sh���y�ؾa�Տס除��+�il0I�a(�����'�Uٌ��+�ѪR3Ϥ4�1D`饴��vB��Jv�� '%8=1iҫ)Y���)V��(�y�`ϋ��X2���b/����`B�g�;��2&.�.3d$L�vL��{F��䕛��	#	��DM��Z��F�����<#-��'{0�q$4pū����3���2Ԡ�HM� �6����e���ʂf}��\e��i���^k�Hw�Ar�c����� *�7� L!�۰]���~�3�o�1��*������
(�����[�F��:�3�J���#}b鯎AҢ.Yu�N݈[A��&��bx���+����<ĤB�H����R��	�A�c	� �6�w��f�.�yVTm	<�����h�/�bw�1���J�}6fn��{B>F,�Ͽ07��z5���N����|'b2��N8h�$&I�nYJ��P�����\M8M��`c�3J��_�⑘�������UIY�z�������XU~�q��t4cY^�����vMT,#'���
V�3�#)8���
�[�kvB'ߘ�����l�}};h��OH��o��6"�пo�Z��;;�w���U���0�.�p���}'���bУ3M���9t��J[���6�կ	C�>�b����SG^X���ɫ�\�̵Sf���&)q�[��MW+�i!E�A�^W~��l�(��Y�|�ʞBc�2N�K�[��]���os>�f6pp(E�f��;z	�
'uSR�:�N|�'���I9p�B�����=@.4��g����+Ӽ4���R�(�; rL��{���$Œi��6�����׎�v�y�=��
:���<I�����U��v=Z�����Ĩ���4�A0�
�c!��@"9u�mZ;�M��z���|�}B�"%���.�u�ޔ��*-+g�3�0���-Er�8�$%hi�r��8[�6��	��b���ڈ���-�[n��l�^m~��S�\��
�)�9p��J�<� À���@%xR�R�]���a�M��
:F5q�w{[�Oi-����x����H��40��ӆ�B�[��OIg��b;WP��W�����n���b��fTP��a�~B���=[z�g�,ñ�����
t�E����j_�<!ع���c�]e��&���d��J]k^����X�]�����f��;I�~��\.gS���+6�nLJ�J�H`��E���Jko6�\E������s��|lo6�ZJ���F�υ�Vk���\r�>���!�zH8?�vAKJ,<¼5'�i���j���~a�j��� �����v z�-����X�l�:�N�fa�p��p�D��f�0\�'�򀸄%g���~M��$����@�V�#|�G�yK�M�m�6�g;�7�Zqq��AmU�6�	j�G��*�}���ܵ����W��?c`�0��^x���&���p)u݉��1���^<)�K�/�D�O�ㅿ�V���CYȫJ�鬏�X��`vi��da��c�;�b���r���U��U��8c�߸�d�A!�	��c���%%s��UBL���4G�����qzӹ�h��T;��n~H���`1Y�¡�OG<���M��h����/ӻf�Y��L5��$@ �o���D?�i��zud�{�j:U��9��2�$]��\�v�KutTT$�QzҽB��t3�S�Tf��0��b!����2M��ǎ8CfCɣ�v�`�im G�5�z6����Af�Hh(W&��M�v�&�{i�����H~�L����Ep���|��*Ɂ8�Z���dH2�R���E£���)�AK7@��Z%>d�O�y�!6a��CY~4��y>9@0�`��@�8������{��h���k>G����yH�q�z� u��4�]2��Fի��ʴ��D1�-n0�x�� ����bu-�\Zbxm�l�p;����P� �ٶĮg� � �
�ݦ���%�2#�ӧ#�W��_ ��8����y��>1߃sJ�H饖ױX�l�N�\���L9�W�?Aj#�ގ�,�/����b�)��\��Q�]��:[�\:��E�v����NL����})t�'�j�j����R'�f������������/�߿t���GI� ͸�*�fq����;�;�؟?��7�-Jn���L�������K��f�j;�ҭ�mWԦ2Z0�ܟkpl+��S�]��9�ww	\��u�(r��y��<�ִ�\��N|�./�
-�$�H����FǅnsĐ��Ow�����k�Hn]/ƹ�,ө��Xb+��#�{N)ձ�y^,R�G�;��n���)b}�(fR_�ɇ��k�%U�[�
�/!�f��-d�����20�)v� 9��1~� �gr�)��ɢ�z4��EA��f��Mp�����7�Qھ{��
DzU���Ul�+���D�?���4��M0���{�$�]ˌ���q�q̏p%-�O�2�ʈ#�?�CN�A���;.�W���g�[��e,?Å��}k���Κ���_����3����D�;�k��I�r�R�.�x���U#��VV����|��P�]���-��F� A���9�j�����dw=�FE}�Ռ�q~��a1n=��ieБ��T;��A/su�0�j�����$�[|O���{���U�%��C�
S�A ֆ�����7Z�N���o�W��0��ٍ��\�O9�SQ�N2�ˣ˿��G��7YЄ`[F��!�=o��	G������j�.#��<��3�����)hs���I9X�Apn�t5߻^�^�AfQ
╫��\�Q��S���m�Y]�pP_u!�P�3Ĵv���Si٫������~�(���4ɻ�6��yi2����N'q&@��E���`/� �8�[Ƅ������r=�w��c%��?X�34,��0���9��Fe��uF�R�]��N�F����V�V`%BPfǀ�n�4�=%����Y��>r%jɏ�!?ѝ^���zΝ�5'6,	��a�l_��˹�8�]f�yc �{�Ӑ��]��){�J�h�[��l��>�B�A�U�\��i��H�~f����A����G4���,9����90�Px�~�3F�B8F�T@>�5w"v
������è¶�ЛqK��������C���K��|wt��n�IR�=��9_�0.�t׿�1����u�=<Z	�D������w��Uֹ��x�ϩ�~�Ũ������Ty���k1���ʕ�i�!/R<�=�0F0��O��!o�2��:����l
�����φ�i�@޺�sϛ����nm�|�{m	E�
�j���� ���nl <+y�/=Dr@)R��f ��k]v� /O#k�m����s���P�4PT�pD^�@,���k�aD���V��\D��`�k�~�V�0�	Y;�0e9d�w���n��>�򮒽\Q3���|('��!��ۑ&Zݳ����1����]�#�t`y���m�PP�%��z�@�KR(+f��r����9&ou�k���Y|���>!��iZ��	u7J�琼��� ��5�h�񼑩�����˚|��CT�)��SZ� �<���p��!4��w���?��g�N�|�_��ś�h9�q8�8]�eT� S��[��O.*L�n`+W^.�.Om<J���8e���<9�b�2#L[���,�=��q�w@���e��b���� ���jTd�[����td��vxc�1ҥj��ҷu��r+�^q�~yo����}���Gk��l���,1��	}ijtXr8���ck%r��#�_|�o9�����P�d�0��Tma���	��֒��N���Z"�6Va�@^�Ԭd+�8��9�B	9�^GD-�V1ft�7� ��F��f���CT_� L,�o��^��=�B�v)	��A!{�"}!ޔZ�g3�9�h��J؉YMF#݈�IP��Mћ��v��ɸ����G3Z��v���cݭIt�]|��(5�c�d�T�x�`z?`��N<˙���a�	M�����q��I�.T\��&�u�X*� �廉VV=�Wi'oLj�S�u�>$�R�n0T��R]�%L�S��ͽ�+c�JD��tֺo��2)LJUD�A:�� @|���i��8U2�|xˍ��2.�ײ�r�n;��(�zVihW����J({�	����ݴ��sV >2�ŵ:&��$_걇4s�H����\�$�Q5�$��Kr��lm �Ҙ��`?_�������?W��_2�l�6a��}a��)'~��@u)��ȥ@\���{�����l�܊F��`�<)e���`��Ԁ��o��²�9�1)��h��0'�0]�oP[�J���:�C���r����!Ҁ0��>1CsJK��&z'��46��c^L�I���J��ô�+�5y}�!ré����7��/�BX��
g�������32��c��V�h�70�����u���i���yU�#P����4;M��*�h�}O+�ejM��&�Ƚ�%.���Fw:�H��U�v��W� I(H���/a�JȎR{�o�U�1m~IS�!�teu��<� U#)Ep���آ��o�����$�0�׉��f��#���J5����eM#c�mͼ�-p�y���4��F!W��o3�����j�M��& #`0!�_�R��S�����D�8�@p������ �����K1�p���a���;4?�|Sl�����l�}��l��@��Y�0��j�ǋ`،��]�騩���C�6{E`�D9��~s�1���e�i�
��&�|����&�M�:�T);1X\
���~8"N~@5O����!�U�ҸW�tH���St}�9�rQ�������U١�������w�B���E�0-r+	U����ZŚ��u���b93��3��u�sam�ב�RN�b��oj�(>�<�is�eT¯�d5��c�aC�O���b�ZP�Gp�z^-�6U/�B�C��d�8�+�ѱ��`�k�K7|�K&rӃiQOB�I��P������v3m�����l�����5��	��qAb�Ü ࡿ����/�mX�h>Q~��2@-čk���)���fr�骀5��$)�e�4iAy�q�V��X5膯XR�F����ig��7�'o�Bk���8!b��k&��u��3/��/�� lnk&޷�2��alK�5��������!]�Р	���r�G�.7����zMܼ�-̨���tR�薷_#�y��WlS�����w���l:��j�&!
��d�#~c�I���8���2	�N)�l�>�ܯ����3�{+��3�᨞�S~�f $�0懊�������@� SRX�vǿ�){R�Ë�\�ؕ,�O����8Ԥ�H�_�[�sn������	Ch��_\S�mWRX�=+ g��&����'�'����1�����?,����6���$��WM~��c��?��<��_~`@NC���0L�T��h���j����|�4�:w��u	�b<��i���_(
���}����\��-ro�R���1-����;X��
�
#R5)j��a��U��W���X��~_2&����˭���H����3�b�w	c���&C!m�Y�3*l� 1K��|p��z����
=�Pmo�A_aȵ�/+n�**�Y�*�-+`~R�v������<·�������L��Bj~�[��"�*�b-�YDo�`gr=�o�z&�Vof���Z�F���8���h24��b�rU`��݉f蒒�xR�������g�<�鱅����b2��/�o�( � ����R�N8�����W��bG3߮(�Iu<a��p'UeD�L�G�YTAE4�.�5
S���F�P�o��$�M��KI�y���ߝ�M���P��gs�aQ\�,&[��#Zs�z֣l�������f٠Rڶ8a��p��s��X��ܲ��#|�����*>5V�<�7B���ähL���\�����$6����&+��e�������ڄ
VT������Sa=�_$^�H�9��֡�.�S�hm-P�ۺ�G��`�y+�(?�`v��U�HR���;.�QO���7��CDɑ�8��p����R#/����m�Q'^x��̌G@�VM�$>��s4v�^���D����؛[��/�&Sv.֝S'0b�I3X�qϾ�3�"AM���FS���Aa/>2|� �!�5/�����	%�	��m�>�_8�����^�=ن���W/p�����44>���3��>Fr�\t=������G�e^���ҧM����V�x����^�@|��8Qf0.p�R�jDNԟk#{�;�#[}�F��nq�n��?9��l���xA�6�$�pEWaL�]G��ib4~_�!0,�#� ҌN�}�i��f$�8���nŢ�^�~l�b�9n��B&yjp�r�
U�O�*�bc����#�}�����<d����EoƺUvsu���������K�D�G�J�6��H���케�`;�_��U)���*T<N;J�K`���S�O��#��P)*P�Gŵ��)L�t�V6��8�;�"2�C� .@op��x��]���w��Z�fR�y�u&��n�u,oFţ���tc;>S�q�r:����8�|�e>����b�	D�R(6��KOjn!pINC2FU&v��Ԇ�d@׎�%��0���x$�a�i�^sSY���V�$#Ix��!H^������.Y�k�Z(}!}�t,��"q?0���� ��F)�����r@k4f�xً�?2+�V��;$�Y{�cO�ɩ�z��ɯn��6��M���x��Ng�A�\�����=t�挸@n��`���k<U&"øP�6mX%�ȍ��P�[+���
],�iRo�sqÎ����k8�@
�N��9�u�M�, �~Ǝ;2@	��d6#��
�{Ǩ�����>䳩/^�h���J��C�/�ɢ��u�����Uc��y�1�H� ���Cڍ�ŧ�T>j���q��$!�y���t�Y��G �/�A��E��\��Q�u�JR�fp.£���1�bp.#��A,� 1�.�� ��.���d�Jc��J��а������1^hd�$�F/����Tb#8�\"a��8�X�Ί�f����=P3�|��]˹��su�f  � �2�7��E�b���xܹd��!�h�ꎅ�7� Q&����j~n�/�g�Ŋ^	X ���� ��F�l�"	�N�5��g�D�`Sy#b�-���,��)��@3f��5=�&�\��cm��6��QH�I�v�x�ָ ���1���3��ߋ����2�D:���x�:���D<	~] � �چ2YK ]��}�`�K݄��7ٌ�Lسu{]��#Y��a��26����M,Iq���bx]��TP�w�\�	:�ひn)(��� ���(�q�6v���߸q��&,�>
y,c^�z�O��K�Z��-�g~��ݢ>���4���7b��0OXj( *��kË�n���L 8�����h�:m[�N�e�{p+_RX�W�����ϕ>X:�Xx�J� BX�9T!T��ݍ���O��A�W�B�e+�����ɻ�%�C�;�Y�C/��d�A��σ`��w6/5�;�N/���B��z�vV�5͉�N<� �8J��#�����V��#i4�瞾��3�ҷ'��h�l�=�2o����m��UN�y+ ߏ������T����������7t�;�)��A���vT=��DF�j�߶�hw��S	N��PQ�Q����!L%���EE���G�bU<����lm./�-rʸ��=��nS������y���a��>q!�l���B;�`p� ʼ��>��c%Ƙ�m	��s +�s5U���	S�J`�|�I�vp��3�A'��-�� ���1�I������Z�9�&H7>z�a<y���f����uf��"�6�\�B�N�}���)90� �JOG�Oi�<�ԥ>�A�K�f�]Q�|�|>�C���C��:C�z#�Y��gv�G�
���!�c�?#1�!C�d�c5rӮD���嵃^����i�~�P�T�b��4��p��JdZ?���0)���A��S�9�1U\ya�H�Ǫ*^�[�a;�)��ѡ���}��v<tN?H�`�~{�_���v]���V��+83.����������'� TG 8�Y+�#Hts
,�lrbs������L�-���^ݫ}��Ϧ�]p� 6N��H3�S��ƅ�Eɵځ�S�G��n�2�!嬑[�/#y�!@��^�(�O~^ o�f���P��R3mykN�E��E^'�Ȏ���D���Y�xt)	�yz����ژ�${����
����{��z`e�Q�����Ά]��2���.��/�#N@�ˁٹe�!��?G�d B�I���DDM�n��w�;8�ŕ=��HZJQ����]9M�t��ib��u"` ���4��jR7�b[-��E�V�ڧs�f�/Q$�Wm�Ɲ0�����������N�>%�8������.g����rm��#cr����+_@�d�J7Y���x��GՒ�`�W�����^����um�vNU{T$�ݲe���bT�lU��^���]i(�=�w4m�ao��J�&�ڗ��IQ3�E!R�ЂeG�e�r���r�2p�v�i_�`��S O����
.¾ĕ팶ke_�Y'G/�*��O�br:b"��*��l n�C>��2i��"[?ū	ys���#v�7�+��vr�s�<��P_���H�^�b/q�"��D�մ��a�^ �?�x����`*q`:����/{��W0�vh�6�x�*za;D($�{��M�B\&�9�� �8B�e��;j�6²�{j���yc$��RE�F��y�&�]�x���h6'����c�RB����e�����	�k[��U*W����i�Xy�˦p����.4ν9<�a<�Nae�����?����3��	������ZX���ł�ZWq�����"��Q}�����E�YT�c���P&��E1�C4S|~|x1}U��7 =>��=���라�N��'p���Dz��|K���h�H�y��J@���4F�;��/��n�"��u!�����v'^�. ��������(������8��0��kPU�B%����0�h����V�m��B��Ww��G�w�p�·�?�b/��H��BK<98���R5�,ŵr�Wo^���EJ�x%'�<��l5�v>Fi��\�/��0Μ���������⨸��o0��2�����.�%Mj���sn��X;4[��o��$������hFW����y�&0C4�?pC�q�=�Y�K�0�Lv/�u!�?xr�V�|� "'�O�-@�������h9]��J�7"ڇ/��pTP�@o����'��\N��c����5�(���d�m���c���`�e�fƠ�A$Ѫ���$�����'#Z��]�	��-�P�vn���j��m�B �U�׷x�"yzG[YK��x��@��61w_������|@��[���z��T�����n0 ��d%��eY�0�W.�{���-n�$��M������
1�Ӎ�7UV�:��zl�1�YS����<�6>1���Z�jW>���B��)P��$(z�&��k3(�$h.��r\PZ�{_�!����U(K�譤b��p<0w��� K-��90IT�Uq`z޵2�Y��P�b����@�'��6���.�4�<�7�c�pb�8�����<qLlW��K8��u�Z��|���LZ����L��[�@����
��5n\���4��M!-#����L�(�TDl��o�S��ZH�T5q�Rv��
�ǐ""�T�D���ed��/�Wg�Z�A�n-��$N�w&C���f�9��W�5��RDU�	�B<ߍ+:čp?�4�a�n�����3�f���˓Z�%nb����`�1�=���ҙP���FMC��:�~�~�[�[��� V���}b��҆�����!�l(����v��ɢ��L>�/�ڤ�<��F1��n�;�h�����F�"1bY�ټ}��}�N��k�":�����'&��fhǻ~�Q�i�O�Ĵ�mc@� @	����ﺳ#�c'���h�)O}������궟��G8`U:���T� �eFH�!=�gh��Ic��"!�-�Q�YWˁ��a����+G����.x@Z*:��p&���
��@�=� T$��2�b/*N�(�(
[�N|1�d_�@D��b�9R���ty���|i�7��K�£�ߺ�J+�}`����H-�,��,�a�N��:c�%���g��w�X�[@��b��?`��屃a15�K	���F>�C�pi�5,D\�N��rA���w�an�w��bɪ�kx��C�^1$�|$�=zEoJ������4����ք���O�:���џ��U1�?���v�#�ȑ����X��ai� M�s}�ǡ��ǚ@N�_���d4n�U�r7���Sf��"?%�!��z��G���4MϏ�+���j	´�����A��M	�T���z|F60	��M�B��ah�::e|x��.�5,Y��*����6���1u��̤��!���P؋�zQE(������8/y���#ʕ��!�7��g�ɾ � ��>�WL�� �H����j�z�)k�U�=�5�Ƀ�IZ�S� ��5��!Q5bW5����)�����&RZ�Ć!�Ȳ��݋�-�����cR��Q١x����ȕ���XPK������l���8�Ϫ�s���Ul>"χ������D��/s���S����:��,uT����=�e��mkW�K"��+���#�2�p|�M�%:�OQJc��@~1��]U�&(#
����\�%m���\�Cv{�l#`8Y{�+���n��T0E|z���j;��>�=��<C�������r�Ex>V�d	��r	!S4�)ͨ���N�7�K���P|My5MHn[��ƾF5�R��ik�M�Aߋ��I��jM��{_�t�g`X��� d�cEyk���܉r�]^�*1��:��p���k���`@�N%� 5��Q�D:��^���nJFB��2f|[��?��ʢ"^�<�q8������7���3ܪ��O�R;@ں���%�,�*�F�E����s��K�^��d7ZF��`v ��0��s��
+��nՊ|ލI~�6����h��X��$"@'	{_^��ưS_2Ѥ�(��s���qx|.��br��L������|T���!}�0�b��t�=�ڤ�c��kC�Mfm��}���T�6�w��}�P����I;z�������d��! O�mH��O>���!��Dp{MA��F&I�t�W<�}[�"}�K&�-R�7 啌�D���܆����q{�B~{�����	�uK���`�A��WA!<q��Z�h�`Rf���u�Y�X��Wږ�x�I���Z�(३���4����{z�Y�k�/���)%;���3�<�!� 
���DP���7!��Jy('�s[{�%�46f�8b��Z]��
�%H�*~�e���g���胮_�CY���fC�ً�RWR���C4|`�Íh�	wOy�b�PT ���c�����s��NӞؠ��h2�䄾��܍�K��,by�T����%z�>��6�0("puTH{�7?ZV�$VܿD!+̣���-w{<~h��.c�C ��z�f Ύ3 ܒ���'t����4Ju�^N۪4�$��mO��<#�&I�9��v���gd^��l1/7Е���	�U)|����*������D�m	r��-9�b�U=�M���v^O���xG0���["���]�6C����p5�Ц^g+�jX�V�!�Q��9Yt��=�9a, *:;@�_=�ibk�`gmX/��Ce���ep���g�>�/���(LL�`G� E��}�h�$����I������	�z�7)N^�|�\�*Y�n�ؾ�/_Ev��t�z'+_
E��]3�W�wm��Rm(?�f�k��t��P�0|�/����~X���}�z'}��7Iǥ1���~a}���f��+$�F�T�J��:p���3��<���\�7����WZ����ԅ�YZ
j ���6$�u���k*)1�X.�ȳ'��4��P�@|��G�B^��B��LT)�,���l���bJ*�-6��'��V����mr��'˄=]�G'I�9��9� �Ɵ��.�b����W��&����GV�Y��3Է�z��ŶzS��tz�Ό����c`�p�o~%kIW�/�k��چ9�,_t���u�=JAi4,�Q���1v�xHb� \�}sr}���F&��G�|��5�`"��*K���Ƙ�!�ߓ�I��>���ෟAC��Y��4��I
k!��6��b&(��Dj�31au,En�����0�����ݹpx	Sڴ���l���(�[BL��k�h�������6U�.�Q�K���'����v��ϾiB��]}(۴i��� QgN��!�aԸ��� �{�"�4�9n�C>"��X�Y�f+�y��Y_q�Gj,���Ű]�X�n��R�+�,Du"W(�2RK���b��z]�<pc�+�y�P�"�u�F界�B�=ǝ5��b@}�z'���Y���A�<K����Ҧłh���ӽ6I�<$�\5��] ;f;O4���IrT�E p��	����xJ�-Ov��jow$�t�:}��|�
X c�1��炲+���w+��A~U.xG{&������*ia+�')i����n�9֍\���ԋ}�U�����͜��H_�Kl��K��85a	�s#u�k-��G�gq�A%����4�7�P�g��b�*��'�j�c�M��Q�|���Tvo�Ԙ�B�g�A*!^nF(�q�����+6�4U*�Ɂ� ����r��Ē�Z�u�V5��%l���-y��h�h|�O��0`*�z�q�O��+���=���o;�\��C:{���0���:��!�:"V`��l��'�
���-��r�u)�F+rt���n	S;�M���*�1�<���fℕz�0}c�M!g���J�t㨛&H��3�$o�,@P{���˂~�i3�g��Ѭ����U��͐N�R�\U��6FU�G���0��Vx�C����f�nb?׺I�m�%��'�%NHY��]��q�y/$����\70g �~},q�{���x���2u-��w����I�0���>7h#)}�qE��}qفb�v�EmVM�ȼ�D{��k>�Ƅ� ��5�{@^����-�0��E�M�YO�J|@�F*�n��8e�K	O�osӍĳ'���L�� �r3T���v������'�y����
��
�aF6����i5X�j�,,�s]SM����D+(��nQ�E�&f^L�"�W4-y�t1�L�k���v��{D��l��Y�lP��}H%q��ۼ������,�#�{g?��x��a�["u�.����}���x�'�h��UXgX��@��!�e���+�~�D6���JP�/��ƍKI����sٌG��,ڤL���qJ���;kݚ��L��?� ��;"~zFD������'b�B֐G�sV���y��xų�s,�{׈Do��<�L	�v��e�zyeUi�q(�v;�:�X
z�`��|}�Ax������an�P��'hp��C#���Z��Vqɭ)��.�Zc
�yε���m�K�W&�<F�G7"j��2�tx��O�O*%�Mc8��i��?���yA{2F< 5�d"��/��_��B�6mDp0:H�Q��ӘCm�hV�+�ą䌤�K\���������j'l��αoX��T{�(��7Rͳ��A�$�v�i��T��:�Ρzi��ZR���p�q�˻g�F�<��o�<�&1�����A�Or��Nd����.i��3���es@�xU�LBA6��gz�A,�	rJ^t��hf�v��n��SJ�9ͰP�aTX�Z`�s�%-~&�, H��f���?���Lh"��H>D���<6����:J��ry�o�4����mغH�/�,�CƗlC[#�ݪ�����d��u}4;��D!�@�u��Y�
����AT�f�x'��3XOʘ�E3�I��j��}P����oRn�?8�5���k.*��}5("�ƁS��G�� �G}M��ր����u��Y��Y~�8v�E��W���q�Tw�����`���BA7/َ�������Π�����z�K.��)ë}�ך�se�����Q6��+,�]ϯ��'k|�#��}<�1�:7�F���<#$��C�,[�O�̈Ru�B��>�a�Xǩ�������4n$���
�~�N��<���~�Ю6��(����ָq��0!��nNe5��:}�ǝ��W��G��L���RF>���=�w�!�h�!PZn?�!���~�F��Đ��o��#�L�{�&�dβ���ո+E��*�s�O�RԿWl*ܴ<ݏE���m}�y�y�\�uذj�<�}�qҭX�R�.e����Xx���xJ���#����h[W���	˓��@�g|n��LIr��� �����T��[���i��#�u�$u5뚘F���@��̛6Zw��֥=@Slck��VN�~&#�����꺎w`:�N��0��g�
�A�v� ޖ�����`���U�N8!���!�<���5�4�C^��KY���Ztz�=�7�q�=�#V�:�זp�D�%�od\[C�;h��Ɔ@I���	����ZᢧD����s��3����E%X�_���ڧ��,�kM��,�F]v�fv߹߬Q84-q^V�~��g�ʻ�|0�v(6��+=L��DL��V��K��e�Gb0����]6�s~3�� ��64�{ߛ��X�m��Mg@QC_���9HIԺ���]��@�(pjE,��C���'�:�O�=hO���'Az�\MI�粨�?ɓN����=���Fْ�U�Zi�H����f{�b��,���'�!�v�F���F5UPBVhZ��U�U_�W�!�\9O��Ƚ����K�c�%����=څ�`N78�
h��yw�������ҍ��ۛ�h�Ɩ�̄������̙�/k��� H��6\��O�l�����ڞ�?�Uf��n+H���f*EPC��=��JX�n
^'n���˵�q�.h�tG���ھ#1ᾰO����\��t���P~�l`�����>ؾ�����߹f>����r�\�$�������R��Q&p���*�D�S̢������du[z��_(&���g�����n0�S�j�Ӕu��>]g�~��\�y7�ߟnOX������C�mi����"��+�sK�,v���o-j��C��D����8y��w�)���kS��^��u����0�"�l����>��$	�Ñ�?�ܩ[$ Զ�l�ۡ^�F��4�j2����|jꆂ��'V]�:􂇓v�.� �T3�5e;@���t�&~�@_�l���
��}�T?ҍ���q|�Am��l7�tS� �#�U8�z�"ẍ�LC��#	�H�ѱ�S;�:
TM��Jc����j>��b�T���zn-A�x*�mf+WM�i���R�^�(��w@��p��� N�;<����c����|��fG��)��-����y}�j�}~kr��T�&��<��|��t�B`�8D^ć���¼�A˄0�"r�^���%���ֺ������1X>>����E����ra�s�g.�ڧI�!�+�9NEƿ���Q��	{����>��q��V͜��{Uc8�M}��p �� m��y���b2h}5K��/f={e��+8i�?��i`���w&8Iö�+�ߏ�ؑ��S�����l=	� ��xR�jE[�y�f:�5ߨ6�DWY������B��)p�������|v�^��	����!��ϖ�ۄ�u�?��!݀ĺA׸��*)�!'����eQW΀�'r��@T������x�%����V�u��]��]����O�H���.U?��j��3�2|��+G�e����a��ʼK�E���2�� �ʹ��:��������?>�5z��B���zPի��_���hTh�d�QV�-�P��p�E���`�'��凄�0�w/6+�?{Ad�)D��'f3��x_�в��#��~^�l���V�*����RME��ӡ�5�1F�.�}c)Ȧ��h���f��0��1˽%a\�����y�R�
Ij����?|����?l��Nmw����(�.�韵���BX'�C�qD�V_��>W�+�AŜ2\�!�N&��(f<��k��`/�,v{�\�7x,T�4���-����-��_�Uvsh��n��?���7uP'���T�?+CacOT�A���:r�#�mdh�ڕ�Ίx��k���W_;����f0N}0�e�}WhP�����BZ�<#�y�z����邳�I+2�s�i` ٬���p����p[{ٷ,r�ע2)��w�6<"E�2�F���PڟT������f��֬�"!&�p5�8�e�d��=�<]G��dJc�����<:/83�ynG�n��vCv�����q���3���W�q�����:�Q��Dx�[J������aE'>[U-��cݏv�K+tW��i��H*P���^��D�D��3�B"��6��׌Ҋ�s�U�S<���c���7k�)Hò](���/�0Q��z�ŒR\������r������ط��5��1z�k�;��7.�H��6��X6"�	���n�ǋ.4�HN8y0jг'�F%ﳪ/�|���h/փJNY4صt����4y;�r3\��a��#��D�4A|֯ح�1b&�zţ1�؝���B+���ܹ�^�F���E�~uX�ΝAJ׳���@�|�n����u,l�2�����aK���K���(-�<����4�_��n����&=�'׳\�ଃ~L�;00�v�-z4�Q5����oPHs�F������z�W��}�{!���h`���d�����P��Oд����iv�w�c���l)�'�=[���ۦ\h��j؜���D3�Pf&�XKpj����,zf����`xM�;�*n�9'�[��S����
�RXd]�׏'��gs��P���翙����{M����n;�g,ߗ��/�mo;��S�xÖ'�8�:�<���+�����@�(t>���zn�X��bb�^�90�w��A�}\�8�z9i�J�0�8�Mu$Q�?"7dz�JX�N!�Wۓ*OU�:�c�lϜ3�R��O�0rչ�F��h�vZB�-�w2�&y�i�LM\�[(a���x���
��D�R�;�{��4��+\��W�,���ɤ��H(�z��:��A�l*tU�3����D��n��9�' )��R*�٤b�K�ճQY۔��'=<��:�0�c��N�4�P���D�-��cNv:	=!A,�HJ���E=닗��mu~�$6gR��q�W�Η�5%�����b�x�ҁ��&��x~��Y�<�����kW��� �����lfzA]#��F�H��}��Wq���"�N��<[��o���Q��m���v�����8�\��-�6ʴ	���a"��K�q��\�<ؽY��߸u�N�r�F�n�\�{�U'�s�̶��ȵ}-Ex���^v�<c�|O�w�u�_��S��n?�u��v{�W�����#D��M��H�L�ڔ�|Nt\�R�h�(��uFd�cz���5�N��|��Ͻ��Tޞt��YP�0��������RN��P7e3�{6b�~]|�Y���d��}� �+X�
�%�`�Nݐ����H�(:q��AR�c=,k�w{��P����yǙ�R�勤�qk��e&iؓ���aB�[u�|E��J�y�K�
�H��?R%%Xqz���=��	=f��:�#���6�S����I��¬�Ӛ�'�
���U�� �n��l*�L�ƇV��A�n�8�qD�WANc7S7Oa�߈Ȩ���#�[��a�/�hd���^��ΒٷD`}.�&;KC6v���2ߌ7��b@�F�'��ֿlb������u}HK}a��{�] �q��3ߜ�x� :>xU�mߋ����F��n6K.� ��P;MT����lZ��.Q����NL��`���mݙ}�7��ὃ�rC�6��;%��u+>R#Ȱ�J_�1ȀZm֪Eވ���@O�^�Ge�`@3�y����"�FF���T���)�88�|k��QQ��҄�)�q�D1��,��<l�T��ٖY06��a�� <��?8���v��/�/�=b�'>P^������>���<vY��q�l�u�I|�(��AA<"����m��J�/��5?���_[��/���@�Tp���Q1�?��H_@?�������nL��ҥH��a������?�P;������c_iעq6,�9����Bq`��Z�\5M����J�?��u��]	�V�C��y�A���κ��Y�>s������_��P+��l�S���&�q 2a�<o[/zIQs��"�"�֕�5��B�K?x�pZ�N�^;\������w�|���h�B"]��Q#d:���6o���a�l��vG	Y�x�b�� �T�+�X�&����cq��M���\�]�}7�؃�)i��R�*;Ͽ��G��R9�8��a�ŷ��xJ�CW�4�o<˵9\�T��Mb$g��(7;��c�:$�k�J��b�P�B����]֗@�fݍ&�x�X�R'7{*�#�Ҹ�*�>܌���c�	kX��S�^�bV�� �#�6�(�sq�����D�d_��@�K-1�C��D�c���6�9�l�q����<j�q����N2&)!O����EN�/��pL�Y@�s�UQ��>.��=�x�����/-W/�%�R��_mS�_n��G{�g���e`� )�ɞ���çn�,�Ӭ�x]e�DPf*ڪ��e��3�rzAB4������WR��gdI�;Q(��ʛ�mB��S�ew�{-��O>���A.PѬ�d�O�,���k�����3B�lfh������'4���qU}*��@�*}
��ߍGػ�&��J���i��_���Ϟ�Y9؀˕�����.X㾲�(�S��o�(L'��V��������,kQM,���
�1���N8�����P��S<�Q-;��vWK�dČ,aua��;�Z�N-0e"l���p��
84uq�9-RlCx�l--u�����y#�A'[�d��c�G���so7Á�0%���z@9mB?ug˷�c��`���Hk%�ūc��ٻ'U���C a��!�1+�[�X�K��Cx��m��4**����IK�%��Q^6�BԌ=+�uԖ���f�I�&B!lCE� ������=������雬4��dt��,�u����K�����u���4��U���v��EBz`˯Dm�fyLd}�Y���L��S�;��������#Lt�Ƈ��E�y_�/+�9%8�Ջ^�x�l�P�_�����P��[5�?�Hd�iG�����o�����
:Ck����
�!@.u�T��)/ ��Vi�7V�Sc]�%�[�(X��ћ<5ۮ������5s���ɘSo��"C�b^SA���P�pX�{Z����V��u���� e����B}��
�����R�w�t�~e��%v����|��6q������ �������??�/F���)e��yO�=A����BI�T���L�cE!��*tqO"�0C6�;L�����WN�ɦ�*��dT��w�s�x.<��¢	VL������(�k?�U��yOY�LU��6���U����6L���I��L�*�����������5��t�]C��ω%���5��u���J�ޥ�r_1����p3.�K��5�<H�öu$1qj���/-^`�<�ox��$�ǿG�nN_�_:�)LL ���E
s"&��g]p�Z�B���nlnK���k4R-w~G��� $�'���U�AG��(�m�OT_�>����Jv�Y�l�Qۂw��>mZ�z��`E��P�d�J4��rI�$D����/�9�Ncg5��L-��u):����?��v
0�����pu��,pM��X��aYRɟ�
��5����&{W[ X��9�@v�G_�tlq� .~�X�}���l����0�ۢs���ޥM��,Ud
��l~<"�c/���ҕKDY���O1}������ }.9n ��{��D����О{��z�Q1%:�[�b����Hv�#.�Dq�}�uq�'�!�N�^�V~+�%�����g31�'������)���կ�PcV��.���N����Y�S��H�|�0���E�����\�u�ׂ"��n0w�����]E5]{��n�F��J����nP�T����8�.��Q
�τ�e8��g�S1��\���� Ӗ�!y�H�D�����y�o�Tl-���#T���*A�=�D>	��&;�s���8��-;�p
D�p�a� $S2-��[U�~���[��Hf%ٙU�/�A;�r��GeV�d<�	�Pa|��:�������Q��q�L��{��N���ۼ��R���)=;Q\�s*2�n���q���|��̧b��8�Kc�H�P�
�`�M})��[p]�����X�}��@���v/H���11=~��	1�����U�㖶�-j0��G����)tW�4ʽ�Z�ˣ������u�/h�R��'�[xF��_�7

X%D��g����k+��m��Qdr�M	���H�kd���T�k12An84)��G.8Sv��|75�'\Ï����%!�I�tf�fa��>�l�mAo��@�O�=x���M���\�������(ڈ�!6:34�.��tJ�X��Gj̃(^1,�(�t����R�&���T��4�c���l���v}������-�6V���>�
�TE:���h��I!�"��ܵ8��K˙*۴��'�ɉ��?�_f*p�s�N��.��u�j�z��ʥec��ц� �\):���$�C�I�%�d���6+1�+ck��{.-1ەN��alJ	f�ЍtaPX�K�'(�ǟBްh�W�mc/�����\�"#�t�"6>���D�JV��Nq?w��I�|��ktl�s����7G�(�T��k@��d�IV��o�!�HP��L�k�s�"�������`0��}�O��@�5R�!Z@=[����]�Պ��To-��w�}Lf�*0�(ۼ�j��)���p[4�tA�e�Q?r=�?�/�O0�ML�f�����S���[ �,�F!�À���]ǌ���+_��t\t/�Z&��Jؿ��P��w����>�R�2����,s�Ck��|��2��z���q
�%i�̟g�#竞�hI�y�4��+H�/�_E����Ñ���*/4��]�o�{��g�x��@�ö�2�sK�w�G�٘��tF�+�hg�c����Ψ��)����72}��pG��L��-���ڑ�!�P��*�*����ǣ̑�q�:���zE=u�y��V("��K��G#>�_y[��.y:H
��Ī��H���h�6e�S�� � F�E����ΖUh�"�91���
�l�P�X�Ĥ�)B�k�C�k���%ӥE����Q�A}�R'���S#��1�Nl�<F�>��;�I\Lϗ���/N��2GF9����l�נ`��:��.�5<,�\��3����ز\̢Gr�`Vy�
�y�lF�e3�g���
�3�܎M8%:Ӱ秎��3��iw$��%3�bo��E̲�i��������?�U,�jօM$|�C$������~!��v��A(�n+֖�=�W;L����4il�mE�L�g����#�b��~��0{5޻�L�QqV{��;��r$��ɀHi�N��G<M�}>�Q��J��]k&��F�e���^f�N>ͯ�š]h�9�>�VێM|z�?S��V7L&А����?ޣ3>�W�o+*��@�N������,&Y�5�J�IT03i2����{)H�m�����ˀ�g��1����#�>$����D�~�h���M�������^�f`X0��V�?��#^���V�E�����{׶���2����ҝ��&��%@���o2[���o��d��T�`�
hC�+�5�MN٦"�c��f�����9�p�wc���-�p��3��w`�:mRt�2V��{��P��kM�����~�nIR��I�2�pO��O� y���(�!�Eߕ��������5��$v�Bal�3��M'�H���gj�*$�2��O*������0��Y��Y�'�NR7���L��tZ��BSNp>�:Yrd��x���P>�����1�ّ� ��o�;�U�Ʃ
|��R.ON���U#t����e>;��l�B�ߠIa��\i��h�V.=v�ĀͼQP;�;�]��N��*#��=�|��6Ҹ����?�!���(�D�z�S�X�xl�����	��ȹC���bGn��̔�c����\A�@o�m+t:��x`g>lw���+vą��p�'�*���kˣ��O��6���Ȥ������]�C(�`��4q�8P�ݠ˕��BkY�D߱��îj�7Ux$0�R	��	�1����	��Q$
�?����+�W�8��(�e�]�
.���؀���k��!1t� �d�g�K��#�^��<�*��U�R� ���N#j�4
��L�Bkr��U"�i�kUҧ���:�~�>!F���-�M����TU�߹��W��T����n��Fll�e]ٞM��8#	�s�b6մ�J�I��&���T̉�!�JtH�ەzh�$��:.8�X� ��k%�櫺�U��%�i׉>�8ջ.uG��y�U���^�ү�ݮ��${�Wj���-gj��Q㌏��Cg����.	<�(�=4_��
��i�Z��ҵwJ?�Y~���G�-�Ƹ�s5���CgR�4��c��a=2��:3����p����|�>d��l���0��F�'3쒰����� 7�yڊ���Ix��5��ϩ����+܋��������g?�%��5�*�ٜ�D�����}���1��&�Y�<*4S�v�6:4�'��!垢1������}����&aMWټ���O�׌~���ȝ��*�]�d���-N\�4�]Ǯ���?�Âp<�b0�rS�P!v�vF��砿���Xw7$�����Ť����=eRBi�>�d��ER���R�X����w�F�"��6A�YȒ����4�A(��K ���Ӥ`�f�fߍf֪
�]�4-����B@MR3�0�_��m���0@�_BA�-GO������&�Q�����nc���,�Y�q~+�#4O@�\.r��VH�tPZ���i�OA{X��s	v�b%�Q��]܇3`�d���]wb����5~���&��2U� ,�(%5�iߤ�-�w:��_5H���r�r�u[/�oT��"�	��4j(��Cm�/���^��R?�H���Ԫ�qr�$��ֻM�#���u�Rj2����wY��_.��<D�e���ga�������]d�����q������~7g�M�D�II+u�~��a1��
	���T��P�#�_A����i��nU�r��َK��Zgx�S�E��~� �:�*e
B����c��k)R�:�7�n��-��yк�ʼ���]�S8b#�a�`�7���U_G�f<�<Z}]�.���!�SI�Y���ڃ54���k1�bz��ǋn�c�b4+�珲�. �[���z۝�d��	\��ݶ���R�_��y���S_]2�&@��98,�	����}r�&58~�=4����͞�hy� 6{&|9T�L�"�ν��r�Qy�|ϤӢ�7+W�!yi�d(M�p%6������d���P`_�	r�"�3im�6����#��T��'(n�����4���\�@��'Q��,�1]p=��(��d�K	n%q�)�D���󱹯s�W����E@�;�tT&��h|k=�Nm�S�$�lX���X� J�e���U�[�"]�7���IY�����G�rZ��u�ݺ7qc8��̊X�tx��Wd���q:C�['膋ł��
,@�J�GwN����������0QSb:�s�PU�����Dۡ ��K���a�e:��|�`rk��I"ux�M�?����~~ƍʳ�I�uu��׭�A5�6�lg�Rf̾c�Dx%&����&V��L���揢�R��޻�Je�6ih򀕮O%��4q�$��vdU�}�v��0�3B�W�J�Y� e�����fv��w��Xg��;W��|d�K|�C��G��k����� ��	`YH���4�eb�3�c�ޗ� s|a�^�����hޖ�3�w��M��OrJc��\�gl��6=hт˜a«g�M��y,rN�H�B��eR�ZY|�=n����JK��"&��`8��c_���+<��"��]䗞8�aʳt$$M*Į2s|����c�Ƹ_���rv�.m��֐B=M�y�z=ʭ�n�9�I��G_5�Q�ԥ�n�=�=k7���ŗ�����xr��c������n��⑷K&�#������F0����� ���n�l����������k�Uɞ�O��CZc�q��`��#��.�LZ��X^�&��M,1���+��y�Dh5搞�.�&�Nz4�5˧��R�*�z�v��`�>��h҃�5��,m�K�嘷�vcSgLzs�
σ�קPYIHz��ٔkS{K��l��{�1s��#�Nz�Twclr�^�-����e�
j}����9��-��9��&���$�Z��_q-=���M��W_��u��oH$�'���r����p�.�P˱�32yL��r^	'�.�Ϊ�v=��t�=rK��Va<?��Y���l�m���[8]����̖3� ��K�%w��"ٚV$naY�ߴ�� t��0����2U��د� �M�����	U5����<Є�zᚸoqÎ�$�MI�l��+Gn��o�CA]U�?�b����7X��]�N~Y�a2Oe�������rC,.1F2����� � EH��yt�`���
]��oռ����OJJK^�<Y�2��)�О�N_//�(�N����;�ٛ�V^aÒ ��g�T���M�>1E1������$���H.o
C�˰T�a
��}���1���~�~b��%��ڷOl�\K�ɱWz�g�FQ_	/�W�	�.�T�x%&S���2��>E��s�s���ٞ��Q8ťO�{�J�Ⱦ��/����9E������c\��7ʢp��W	&*�?-Ŝ6	�i��
`JA�y�i�fLU�ut���,�5-��(�!��g�k���L�ʗ�;�u�[�w���lX�ģr��3p� �?��11��Y����v���os0l�Rr�_������ۂ�UæBE��p�;�����eLQ;AV"�����]_��8vm���i�G߁N�6�#��f�}��	�#�B���vf�w�|�
���1֭	v�<��୏�m��:^�[��d�o���B���c�[F�MO����J0�\��A�/io�=Rvw�]8�a��א��܏j^Cb">!��D�e}�i]Ժf����G��������".�Pމ����'�'w��o�Ă>�M"Ɏ�U��2�+ʬ����7L���eԭ/�P�O˸���K��v'��z\��j�.�?��f����o��O�=��H�K�c�m�5D/��~]�!Iyz��՗-ڃ�Y����n�f�ƢbH�؝���T	?�x�U��"{���82Je� d,`�m�q�w5n4n#'=�^O��wt���W��}3U��~����<���HY�Tt�O�T�앜��pZ�CZw!P�-�br��&�w�f�0Up�k���Ζ�q�rW���
'=�<�1�\��~i������:n�UNn�۫���\�����}��Z��xT��Y��w��Ak1�����pLwN�@O2)0\3�jA�����<��o��żm �o�w�V'���j_�o*V�u�>�Km����Vn^N�# ����8sE2zr�DN�����8B~:W�J��V�:3�d�Qj�K�^�f,:�ˉ ne��ƿ4�7����������O't~�R��xSF8�il�$:N;!�bʔ�f�m�W�~�9NP��V
����0�7!u� �P��h/j��xSUSe��I�s����f����q�@�Y�H��(4�h:?U�q�%�c��m�{��9�̙ubBmyl��f�+؉��s5��ēF��J����:�^r��|�ԓ���U�x�AGEtJT���Ӷ�}�
�V:�ArW�%v�P���F����>HZ#�d��,h
CJ��$��D�����<Y��*~�"��'?��°D�a}9Q~��\)���Ͻ'�t��n�z�5��rkU)�V+ ��������op��4�-��D�?��5t؟ ��ÜZ\ �7�˜^�}���<��UM�:�>���+��K���'S�3 ��A_G^%��uE�^��cX�9^�	�J��屌���$�5���!�r�Z�M� ���tɵ��H�7n�v�38�������Q�_��b3����.�<0ݼ!vű��|���G7�UhR�1�nO��j�8q�G�1�N��
᣸�K���8vn����a�{�@g��F�l4�#�x�d�`N�tl�Ǟ�؋� ��DÁ�Ȋ�1W�'rh�T�� ^xT8�z2��.;6��&�
������E3�FiE���C�&�zs���k�d8	."���wY�C
εMƤ�תdx��{��t:!{O̯Vdr�J�(��;FZ�T�����o�o=��Q�̯^'T���P@0?�o����X}��;4��'d�?��aB0���V�qs���%�=	(�������e����Bv�0���5�R����L�y]���d��o��o��~K�s���i���;�R��xY7�j��c`C������Q/����������m��rRó��l���U�CWIˈ�L6[�!РnD���Y���yTq����Ȳ���z�mR߂�w��i�I=2g�݅�`���G�X ;��<�+i�?�'��"�w-���k��yȳ28('�`ܫ�����{����/��1�J@�+��?n�pnLLjȿ�����( ΅VX�tQɯ���jû��\Т%+tn���@���i���#D��x����/9I�XM�ۨz^ћ��!��s
�bѰ����`�EdRD����wS����0�kԽ�s_�r(i,���N׸�d�v#UD��!�&��|���I��+�U����ˣ̳�TE�P%�f2�vG��L�]� �f��v`��sg�.��=�P������<���G���^�4�ebx0w� #�~���1/� I1�� �w��y�����Z��E���H-��{�bPy烦	?j,D��?�u�Ea��/Z#1�9z=���|��C���g�O�ET��y�X�$&cd��b9�CA��^��%_,�{2}�rX>\͘3��mY�g81h~�*C�O�{�N���>��d944G>O�v�Qfi*6�K7�a|���\I[��a!<��o����%�:�~�]�vX�,s��E���L� �~����2�n"�U��<�xE��ڏ�@���w !X:&$��=�
�|�Uɫ���d:�*�/�ܱ����>�,̏��08B�����[�k	Q�=;ŀm�#>���������dge�j�ń�c���2A8���U��Sz���v�A�O�}�e��
v�R梌�����'aݺ>�&`0�mä &�kZ�"�1trǳ>F������2R��� �\B�
�ӝ`�C�'���>����r��+w㹃N�>h�[�v�U�Gc���>��5rN�Un@�\�/Yt'�_����ZB�Cd��r�q�@߽iM�>��/>y�����I����-˝ǉ�̡=��{���V��]��b�ܨ�ѿ����]�����(l�8��������Y
}��Nt^� �;u6㹗��_���aU�P���dp��Ǻ����]@A�Y%��d�Lo�:_��i]�淨��Y�>�Za�M�*�h#)ο,���O6<�#W]�Ԑ�qt0XD#� }Nr:����-$,�,�}F��F�Ϫ�Z�z��gf,+� �%]Z$j������i�#��ݪ��7��Du�v�p��Dy�ESN�N;�eR9��4C-+�1Dz���ql��ӂ�͗T�ٯ����_y��$\;5 ��}��Zǃ��0�k�Q_�s{�U��N�vz��@�-�т���1/�V	������T�zQ�]eJ�lRi�"��ޗq��*�^E{��2(��|\���hJA�����A[���W�&�ސ�:h�R�Y�s�H
%���~=�C[��qs���a���w�5]f~�bl:-^ߺe@Wd�?Ё�c�K�<�v�:ݺV�k����cۉ��� 5�k���� ��p��J��c+��Na�k��+�i�Z��nF�1(���a�́�YD��"�]�s�J��y����������99Udtb��Ϲ{%RNBmE���<��:�Vu��̷�Q��A
0�t[������Ig�GW����W]߈W��r����$<ã;�+�}
��Rbo�YzWi^�O>�b�v<��	4�%��T�$4�?�����Ќl�}�	�،��������j��в�Y.��Д=;�vwG��?�# CRy"P �n���·�A�Hܽs���JfDq\Cj�\�1�萘yI�XJW�L�"3�
�_L�gRp\-4qR��v��H�P��#�(��oTeiȤf8���8���}	ob����[VoY��<���
���AQ�J��ٺ���,�	ߑ�����@w��tW��]�N���{��`[���4��=�AfFShD�2���hqL;��ו@����UMiS����"��,��Y�W �I���Dh��s<,����3f���D�n�nB�^�B� /쳎jBBD�+
Xx9T��t�t~����e_��67�9��/�)�?N�Ȉa��~0F���WXە��8`qn�΁t�!���w�VɬΨ'�+��Y�1Z���.���&~Č��S�Wg�$D���+7`�L��w�Ko�O�OW9�QrB�>���D1}'f����U��l�ʥ-r�i>��j��)?2��E]/����"[{��Z#.��uv�Ww��Y�A�=Z尛��EǬ��2~#Jq�d��f����z��H	�D�;�F4�2tL%"ЦB���� ���T�������X;�GP�{�db�@%�Na7p��0�.��s>�S�3�
�76�Z�6����L^��r�id`�ǢA��|B̓�ؗ�~6��(�'���Ri��������}}�;�%���|�P��8���ʑ�/�+%�Cl��<]��-�]�9q�ikY��qHVUM�H��j���|֤>cM2̆�
=��7���.j[$��Q$� e,���!�p��4~A�b��C������ve�����3q�����l�mp�H����>�[�������	�ďiV����%�.��v��]<��ƭ����h��c3��s��ݶ��t��,y��)�}�\���-� ��=��1�V�f�9��&�QW�%��n�]� ��)�ās �	���F�=МɲQ��F%�U7���yI����$���ۅ��Z�����U������]"���]@�j������~��y�H�C�vFٌ3���"��;��rwغ� �d��v���m�<��#��n������s�Lf�j�{L
����ȑ+Uw Jd6%$�!��PM)�p�\�^{~���_����4�Y	<��p�]J���#fm�+҂�����מt �Dl5��]y�$��)�ż��3V8�j6�<~}����*��@^r�p������
��h��Xĩ�8�+��M�:3O�`���W*�*�?�C*��]>�S��+	R�s.��bf�i�`�,5�;�f�16�X�K��7��#=	��@���Xܘ`��L�w}�^r5�0���������nu�>�|�)-6q�4[�^���j��%�36>�km���4�(�F  ��3�u�+�2�m�(��(;��������2~��GE��L�s@��y�0o��R�,З�'L�O�h:/0
��˱���tw]�0q��5D{� �U3s������)�e�Ow��Mh1� �����[g}��x�v��pLWKKS�{u�^�Q?��%���,ެ���4�I%�.��fS�2#ꠕiKCF���p�$�r&�'�N��d��A��ף(�����8^�9�?o/4���p�N^���'��:�d�u�r��������� >/�w���ǎ���t�� C�n� ve���K�Q����G��u�Ҧfv�f�8���L#�)��%�}��PQ�LZ��]���,.�u���@�gW��z�L����,jL��T%�S}��k���)2r4�Ǟد�l�	}����fqk+�)�*``��Ma͟Kk�t�Z�Rf��/�m��bc?�ښ9H�ŏ3��k�)X Y�f qN��Q�!��Z�1j:��5��UFD��J��&A��")�rԩ 2����)��!��ԛ��,7�T_�f�Ԑ�Z!�|��Gu�v���C�p'H?�V�B'Jm$�D/���߅�'�D��TZY��?s`БFՑ��U�����w��ș�ĪH}�ѱ]*���M
��n��9P��Z��}I!^"�+�f�Y�	`"��^�w�f�vl�4	n�)9��h�~ù����G�$�Y��^)�3<-�8���{��w��h&��pO��E)I~��R����Ť����EO�,0{#pĜ�
��)ʹJ��!7G�B���?��9[��"O.$M���DfQwA6G���z��؀:	1<����զ*�,�"��O���67ma{كF��0�V(��7��'R�����?�P#�_�n�$�&��S9��e11}�%_��r���l���r���
��g��=3,�qZ��)�r�q;ĳ�y��H{Q��!CY�6�cfd����xD��N�H�^��9"�n�,D�p��O�b�jw�[��c,S�]�0���C�lD��1��{��1قD�T5ūa`c��,
�,r���w�浓b�N��)�>�������l���,�C]!� �8���]��%�zc�U�-����K?P�j�ŮxL:0|�֒9>�;��dւ�&�D���[�۲z�l����m��b�����\B�	�[�.����w,�;���m�� Z� a�8D3��s�]����>�E^�3�$A��΃�O�C)!x�Iw�B!X��=y�Q]:�N����^p������A�TJt��(�Q��ĳ�fM�y�^EW��{���P�%����/z��@��֪Qؖ+s�ʐ�	�%�x�]�@י@�6�������$ޯ^�+�vm�	��m���+��V��`��tۆI��J`Lel��(	|��_��� ��5��GY����a'����W��V����!���;���C^���J��V�?�&`-�sD�F���*�'�+T�=n�2k)��=���e1��c�]��@�6��l�0�
�I0y³�I�X�3|��v2���9D\��s�Rm�σS��nP�c���M\��Wp���I��Μ�������}����|��C� T��`���|�=$u����k��ˇwi���v���Ha�Ke�u���Y��/	���G�N�s%W�P�<��B~o�ȡށRЯ����$�p�Y5	q�1��x*���ה�`��CĄ�������^�C�ˌ�%26���,��\J8I��T�S�^�p�%�1ϯuǥ3���}�HlA{Sږ�����C�>uZu��PI�щ����m�T�L�&��qB�{& ��V� ��/'2� �A�s�;�6E
v� �RKF�E�I���ٵDU�������ڟb+z����Ԁ��ŭ�\�2TF�����e�6�l�pO�J{� ��0��TD�ӄ������A�̨<�"o
s�IF�U�:���}H�����P���-oO�L��!�r�	*��q4�d�������̊ˤ�Q���O�Y~K�G,>8� OkX�����s}�1��o��>�<*KM���	�ϑ�G%>T���-_0�ծ�h|�x�T�&�����8�k���+���g{ม�b�X$���.N�F�M �U�B�3���)f2Q��.x���B�v�� ��3W�g��<[�������}6����*�}%���0�����|&:� #&70�aϛg��<�ß�>ѥ�����(D�o��,]ݷɐ��# �`g���y�lsԈ�x-Z%ќy^������>g�/��m�3i�#޾�;%3zt�|;]���x���Ȉog��.n5\�%*��	n c����%�$�5��v�zy*P�&2�P*��ټ��ǗЧjX���^0�\/H�|�S�>�;�I��E0���̔�v�Z���ůZ��]���ƙ��YfZ�� @b����9��$�k�4�g8IO�$r���,0��Gd����T���@�τ	��J�"����jM��%��ȯr�
��]Ywς+vz�% o��`��a<����U�U��ۦ\oe@xQҶ7��a5���Ͷ�K�_~*�Kl�V�mD�8O����û�cҌ�k־�Nr��Ξ �mU���B�������Vm���v����px���\ˀ.;���^�ZA�6Kv��E�э������^���"��6���*��O0��(c�>1A�(�
ȂqA �!��h ���O�	�.i���O�=�c�x@�L���Jѝ�CۏTyp���lK�B=��ja�H+�3�JŴi)�%�i��=�ZgHTEYd�#�՛���=r�l����I�Ի�\���*���F��R-*��QI�ﾹ!���=Ѡ��P���{�����*+Wx��}&�&!/C[m�Y*ّT�M���k���o�@YEra������7MET�X�Lj�d S�ef((pR� L?,`��t��aG/��膋��X8E�!480��"�>�˦i�Կu:7U����^IT77��E��4i%�;&hE<���g^�W�󗭢s��F^[-<=��������r�\��(�Xl�G�2��0|c�_P�'���7%湌�ǃ�`� %D��ﭻh������Q�eH�����?B�Ue[ U���)h���G����0��)+��9oˈ)T�<�w{ �����YZn��y/��h@�&:p>f�5hA�kU�e� L��ˍ�o].ͲH8Rp�#���{\�7Ν��~+��eG�I����uE��c���5��~Or	���������e���9':��{��4S�#�q�\�pl=[q���ih��+?Yp��aQĂ�3L��yVq�-�W����t���n3RD��B���|>).y�Z��2���K[����&��A�>�"Z�C@�[��vȓ�� �Lgd���5#�KpMr�z���r�b����/	�ӎڽP@ؒ�z�Q6w�z�x#`cu	ԓ~����*ot�X\z�+�q�^�4����Y}�J#�dҴ~�fq�����
NL�V�	s���l���לwg ���2���כ�r�"�٢��&�/fG�߃	�DD'CB �ǀ��։9 _�09��lo�nxN�[���B+��R\�&��%w���僛=���Xh!�P{
���Y)ź�S������ΜUzl�R_!����yYN.��T��yu�O�'r#�b��J#��TM)���"d0Bw3�]��o��(cEl�<|<^���T_H��E�o��?���WLf�1f;��U��N}P�*k���J�����F�m~�N�� ?q���J}+W�Ux��H�-G��E�^��_��Z����''�8������4��Z	�T�ݡvt6����_��b��4�^��Nf@#�#���ǀ�1U�n6�R��� KXUtUAQ�r,��ts(}1��i�����=�?g��)��4�.r���_�P�n��>�G�l�� ��Md�͂�3�6�3��DB�1�C #�;g�!��˨���?���`�0ɠVS;�EE!��*��S<�Ù��,��V-��?p����
�>c���)���[��I,-��F�j�y��STf��t�K��wI%vhn���9�)�1+���pD�����z�W���}#�>Z@c��2�4!{&��)�p�za_a��˃��Ϳh�6e����8�����3� ���?C��l�P��Y�@?��p��"�u�=����O��������L�/��$��L���\����k��39�|�1:dYw>E<�����u<�V�����I�uy3
+Mu�v3���T^�H�U�C�;OK.h�7��W&O�Q�Bh����>^�������+�T���g_=��$a�<*��6��}�Hh��J'4i/bK#�2�Ij�T�g�BF����j\UP�l0��_\r+T��;b����%�b���%t,�P��v��iY�̏(4���`g���3������I�qc���|h�ٜU�K-WADz팰CxZP�L�~o����a�XD��(��_}���=�#U�Kk��"���#=�~�2�D��l���>�����;o.�f�;�Q�O1�-�����,^�0�B�fc}�Y�����3W�P�h`�M�[v�O�!�1�H�z˙�#�ذ�=��SP%u��}���a��Y&>G	fO,�I��â���Qc �%_[Y�^��2Ѱj�0�����&ET�o8����u.' 9;��d�Ǭ�^�s��ȈW�]`�K%�rg��ϖ�RZn�z���S��cH�� 4�$����VioN�P���mX�u�}�|�g�cJu�\;؛��=]I!��|k�#x�op������F#�9p�.����j"��hK��}7�~�F�.$P�������~��jHs�6�j;
�ն��:�;���[����o�)N����$�Sn�C�7��:�/T-m�Tl
���I[��y��?��OF���4���م����?��mC�C�(y���:w?��������f�ޅ�x�ϳ����$�|"iX�D���̝-�+z������E�~_�s�ԡh�@ ����=�H�Ojc	�|��";�{M����ڛ�X]�9	(�	�������?U�ʀ�ƣ`���p���%�#a��a���c�z7jw���O#��Ő�,�e�ܦǭk�<����r�2x�;�K�V9�y����+Va��V}�K8��|�r�㱺��?�Fd0@1��!0�4�?�c�z|YH������x���� Yk�$�y��~4��w��LZ���E�Ӆ�˸��r��c3�g�7���z���֐b�����x���(�6>1� �<	��73��+<�XQ�r�DA��0e��a-���y�N�.�#됮�8]���X��G�� ���CEҴ�7	��-���w].=p�t��?�/�Ω&�q�"Q=n<k���ⵯ�ޠJ�O_�RT`﫾��$|��$y=eS(�q+2������P�r~a�ү<�ߴo�
��\k�$#�t-feP�nSM�t7�BQ#�s�>��29{�����{�l"n:vU��*ps�i��nU���"�	��s�1���K!3����C�/��p���v��"N�Lw2�l�(��W.�sa����ӝX�m,e
�i�|	�͂�oL���H��-�U�.�I��;<��R�$�f��[�4�(�To'�i-�Ľځ�3�Z2�M���]����%���9�Jľ?@׊�]�*��C(IL/ҝ��'p�w�g�b�ʼ��>}҇��[dm�vC�O�W�3��w"}6ё�L���Z�B�ӞƷ���q��f2/T��
��3{7�_A�\ͳ�a�W��Bǋ� ��7'GVh�Q2h��i��km��θr
���@.r*�b1/`i5;��Nv�۴:�d�Ϊ�8 ng�KC��RXHj�=h���%������&/�CO����c�����[����7D��B
�"���M~����.��|���'?���<j��%��E7�PR�۾��&%��}���;%~�d7��=�I�~��1�`SS��v(���<n8�z���D.�]���xO��T:���X��Keϖ��C����B4�����'�n�ʨoC��]�-��5����ڍ(���s&~Q�v�7	8
l��6�h�}���CĪ�;{\��>e�,��|���%�z��u�	����y^2��7|��;Z�T8(4H �;��<��6�Y��g#�s���8r�m4|��i1N���E
�����c�Bn����X�)�`I���1,�y��tl��l9�� P�W�#��ij�X�� �f�Le �i���0q��5+Z���)��3=ҩ��������pK+��owgY��mG}�o�NNE����Ti.�F��~�����'foER/?��_r��~M/}�ߑ���^���7C�G�ұ�_�W�����^JQ��5���?����o�r�\AN���d�&���~�&Cul}G�(�o:�3�Y�~�~�(YrL�xbd�\���T�I�O��#$�i-�lߺ�sUhv숸aݝ�F��#���NU��x0��8C�n�:=�)�n#��nk�y&�$C���A{#I0�/O����D}�Y�d.�t[��+�/�>|��I�p��b���Gy�}�S�����X�
���Pp�1yZU�E�� 	�+�iwyՍ�:� ����vB6�o�Hڹ�Ğ=����މo'���ѫ�2�1q%���Ǳ��t�!w(�Ҭ��by��O �|�R$cH3l�<@��g��|U6(c��d'XP2�l�j!	�p�Csb�j�IY� F�n��z� �U��-�m��=�NxN3o�x\Bṡa��x��O}hT�l	������P�m��5����5��Kp��4�:G�fJ�"�� �vB�1�.�唎>���>�S�,U@��@UE/��6i�*����L˷���gJ^jC�NY��?�n��~�XfI�]��v翆���$�+�<I��f�.��
dR������32�2q�����a��q~g���.���;�?D㏪�mO�0Gj*A.y�<ٖA!�{"=�n��&LѰk��;�[��:�U�U�档�a��N�,j��@�=OA�>\����M.��7��Z�'N�*N
����O&^vG�/�����ٰ*[�n4���H1-2S�ua��lf�]�G{s���g��v��>��X8? ��x��
j(>��q��ϡ�r��n�F�4&}��{�Α� )-2�s�;�-2Q���c�����L����\�U�P�:���]�Y�"�����	;�Ŕ��E�Z�������Q��6pM�"�)���`?�� 﨑C�O2�V���-,�1y8ޱ�>Υ��m�V�0��f�=���]��'u�~ѯ/���8e�yp>�\~U�-l�qd�2�T��i�+��軉#ͳ��f��i��U͗V)�۰E,Hw��m@]���K������Ni�z�,��]��3�e	�)���>�@8E�(�����3{ĕ_핎�������}3{���榪TEa� ]r���	Y�$�����I�N	lu�md�>�@���71�~D�e���¯�X̏F4�N��;)-�+�6���i`�-~W#��r�N�Nk�>t39�l���{E;���a�9�r%�d"�q�t�+M=��Nc�0�鬬j����f��>6wџ�Aad�V�"M5�\f7� �V�F<��p	�NǢ�ȩ�����Z��h�GS��_n�7�y�y��Rۅp��d>��4�b�eaD��(`{G��J�ZH^R�@�$�����O/P����xE'� �\�p�O��j����%j�_��-d�)m��S�[�;����������QW1�N���l��G��[�q-Iۘ�N�ڏ���4�z���ϛ�N�����0�#�|5�a�S���|3���Px�f��#Ж��2P]o2���u4��j�0C������*�2ǔl��V�5hP���e���~J�=�KB9[�o}�b]U�x�v4�w��˖�8Ԉ��Ƅ"���q-�>�f�F��ۮ�Da�\E�0�"���3xi�E�	�|H���=VR���<��d��C�S�d
������ZǨ�Bj�W蚟G^h?Ӱ�("e-\�RU�~-�"e�g��N��3|!ti����A�	��#v̂ gae�
-�㒼���7��U���Y}�>?P/��T	b�ܮ��}a��A�9�~i�wueN?�~�LsIt��7�7�	���p�	`��_�l�Uo���\��_ɧ�A�����(�S̃<p�6�ܺ1V)忬W�̝��.�r}�$���n�K�\��/ɤ�=z����/���ice.�3����$K���ѯ��<�����K"�5�|wAܦ������t߬\����.Փ����+�zW��kc�5��W!ٌ�3(��##c�f��Ȇ`�35���t�(���z�{���p6�r�&:;�^�<�qnv�����7�8g;�2�����'�ɴ���I�c��Ёd��xr�D�h!���c�UK������u"SE��<�9�A��H��Iƌ�@�� eiz�{	#����wٙ�T��/^��k'ZFgoޝ�]AJ�ɧ�N����z��~��&��tGj&N{Kt�/�M`�3X�l�c�Ly]�~�d�s�R|�"t.���$��;|����V``��Spj�]~<��=��t9����q<`v�S�a�W܉��E<�='1Mìzs��Zp��	����Z)���(��lc��z�Sq�Y�8��:���F��-�}�p-n��m-8��XP��6�y�L�]�l�+PŮ��$ l .� ],�j�85�bOA�*Q�a�2��Q�HNf�U�B�_i� �a��f��A���3���DHC��9�]�.�w 1�xmD"�v L	 =�����E*�B�,�L�\4��4�b2<�sй��a���K���˝�s�D���Z\7�� bi=;����t8@V�LW���I�ǃ���Q�	��Pu���F��@%'��H����>�-�Ө�r�-����ɓ�m�pbKQ��>صU%�I��q(����=A�"T_�U������M5�B�ac��쟥�q�^^G��3��'���P�����p�AN#;z|}Yr�� �|R��)�Fj6vyS�p��>Yg�<��=���V]���]	}36�����E2����;m��b���mH�U֕ƾ/Я�O���1ȨC���\ �Y\��V����u�N�Qۓ]vs\���خ�z�=�0�X���1v�|���~fP�.�!,?VBt�9;3,��"S/X곑�2��F�f9�(��?}4��g�
��t1q��(*<��_���	���:�	[���Fl�c���E-?�v �MvY�P��L�J�ٹ6�XbJ3|�>mi��gK`\h�٢�K.��v���0���������~��X�ܵ�L�0�{UNs��'.���0���m���H�q;DN���T��+]Z׸�)�Rr
8�Morr������lllf�%�8i�n�/4�T��K��]��&K��Z_������5[s�'�%��U�1U��
�C�m��_g|KN[�y�z�TLvƲ=t(0�x��0��t�}�fn���E��<	퍥X�6W��q%a%i�Z��$���F��8��IVU�,��K,����%���G�.��F �|��ʫ���Z���[�F��آ�����E��?��]�-����Y�M$���Rz^��m�*!�kv����%T�z�U��ߕ3�z�E��^����5��c��I8��U����)A%��������f&��Ę�iЏ�P�P�a��\O�fF�����J�e/L&"���\�ؑLb��(�Eh����N�D'F������X�u/�Q�I�$}KV"�X����q�&�CN&�.�2ʰ֎�B� �:Ն���#��
��#eH� Um������P�/0GE8����/�%6sI.�,�բC,3�/a�;h
�&]Hf����u�����lſ��]���O�5�(�qt��C T�]+,�x�������ӫ8�h١�±��me�I����sFۜ��dS��[�.���Kli�g�?�����aR$j�h��Ŀ�2ˇ��p�����R��d)��������j���x��d8V��Jv�b�k+�%�Vb������ΌG�G�te7� �<�;kצ�N�3��"��)o}#��o��C�_��ސ�|�öL������:� �֮�N�.�І�ئ��&�Ӵ\ vG;�3 #�
��y-
����|�
<ߗS�c��+F��4�!+�]h��r9����I��G�A8�b���1M��}a�|��s@��c�(��9xx9�l�K��0��:��>�Q[�yU���/�	MR��.�!u��=AKP��ُG5��؉�*�'4��t;�,Jy�\�O�:�8c/E�L*B�51|��R˸�e�H�FİY��|� xv;v������a��Bi�@�ba�����x�����/[�'�,���Gsc1���w%>�OѶ Ы��-�RdN$8��O��9da��<a
�ь�b�a-�=lU��[!��h'�v�&���bg(�C�n�ذ�4�|���q^hʬ�W�|�j�FX*�k���i����>}��N�d[nk�s�EH�	Ë��VEq���g�,Q�������U�Z�.*o{@h~�}��a{�·O��I���@�L��é6�U/IqbQgF_1���5J+��.J�U�״�9��Þ�*o�����"�Y�S'����'�C���lZOȜ��\�O@S���<��i˽s9eUV�z��g�X�'6�a��B���&�j�=-�{-����w�� ��D�o
�cL�Z<w��1��Z�X��·���@�-���p���^vRB���s���:0�oȂ����)Q �V�$6kQR4.�R��>h�D��ʼ��V�q��L�5ZEҬ��Q�p#���NRR��.ޢ11�.tB�Ϛ̦�$�ӗ����{]��<�ɻS�;�dy��&��\��L�@KK����[M*7�h�?�`��7B���TC�I'c��{�ݙ��l+�Ej�[g��\�(�dg��`��4��/!�v >"����r��ݭ�(/��ݧ��� ?�����<o�#�U���[T��ƺ�^K6���/g{VP9�Bj*OW8D�Wx?nd��!�9Y%�g����$5λD_̰T1yb������=��(��15�|�,��jPr޲Z����Y�A�b�fHrGQ�f������2=�\.�W��'#���:B��a���D�lew|Y�{-��LY���Q��)ZRo
'W%�3,�sN(��q_y'9�R�uf�l�7��l$��5�"F��-��d��njZF�$���� }o��b��Đ�'o��9L��J&^i���c�ld?婜�<���ŽN�T�������f������9}«8�,6��8��9r�GZ�ֱ���e�N���xDzyG����@yZ������f#��K,C�?�ivՄ�*����4�.X4��[��a�a���`�4׿v(	�c�jJ��4�Hv��W���Y�(�o�g =_�si�B}+&��`�K��ʰ�Y��F����@×��D�wv޸������o�VO�Rw��(RZzPX 5���?�K��`q�l`Bq���	���J����S�j�L�H�?�����W�aA1�m]�oVv���& U���"%�\F��<òJƐ��p����%t�9��q$�g�NXlf�i�L��oy}�F�j1l//��w�5h21k-6S1��WTe�&1�����5vZ����:��ʈ��E:�����Fj/�����x��j;��E(P���?��,�!ѐ�%��*���P���8%1�!sl������z���0�{=Ȓu~`KZ��$��&�M�A���l��h_��Xė	���iQ�wL��\(�Ԏ�}�8\�5��0c�4p�������^�;��hS��@��	E)W�	��ĵ7;�������K[�E��$���V��N�ut>S%��T\�*)�<?�<&&��`���D��G�X1J��v���� ��;��&��?N�D+���g9�`�Lb��d; �I����I[��*~�=@f`��eB;̦��<�d��rZ�˨}�'����,������l׀HL�����ȑ�;�������2{PGTk�ڷ��Lڛ���"jP��چ�gD��)Jׇ���"b&���ќ�2�Kp\��*я|�����e>b�
������ �U�����݆�����I���`M���Ţ
���dL�'��q���B*Za�ȍE$����
F_��N+�i���\|>c/�P`�mw[WH2OKh���D+�М�Y�Ƭ~��RHNyG1Z�Mχ��Ƹ��I�M�[i YF9G)]R]1aİ��~"UE��>]6I4�Gy�������]��O��h���Y��R-!�t�c�,��X7�4z2㴁���mԶaS���d��
�����	�d�[���n�q�c:bB�L�{���N��6()hldD�BgM�)�OFb�x�`�x��;w
Ԑ-��"��������d��9������L!���՟3����J|�`�IA`D�"�N����t>�#,��E)' O�����{�k�0``��Fxr��شoGb(���}�� �������Ǩ[y�7D땺��ō�}]�0@z��}�J�
��	.�.A��'�9�C�fhήG�Bw7�X��m"���g��kVX[қ�6V�����.IM!]��O#f��t)?�ă����«�Uب�G��l�wpF�u��e���ګ�}֏��"�&rr�4�E��9n?Ox���:��M7�6r��$�L8��'.��\���+?^�F���
�.|d�;�>ó0�\ 
f ��(�}��+���ĭ���I��乙H�w���{�ʟ��-�Un��o�v��J���	�3J��l���9g���kw�Mm�U#T��o@����nA<�N�革*C����p�{�]̱�EJ3��w��E$���PL:}qdR��-:&j~��KN/=�1�$���,a��%��|�]-}��$ڂQ�K�l�e���@��ƚ��P��K�����bj%Ղ�Uț���[L��y�!���U։���c�A+�C�r��������\����$��k��W�@�3�N��$:�A��h*h/�lQ��s�B(�g� ��W�=����ޒٛ�t��F�E��p��-������ĆTo㊴J������Q�~H�m��cc7�D��4����I�csL��!^���9>�J��/D��,�v�ل�ʅ� D��ޅ3��/�ؿ�[�^�q@����zP��Pcj���n�}ViG7ʗj��$Q���76����g�N���~Nπ͋/iU1E��Ş~φq��8
K��b%M�CE!��b��"�L��
�P����5E�Gҥ|�R��o�c4��Jw?�xZ�ǻ�m)�ؗ�s��l�pqX�O�Q�&s�ׁ<<ENi�%�Х1Q�t�u}�+���9�wyv�_�-�V'�C��O�fً�:/�l���8f��Cy�mȒ7Kqc�.�+(�'ٯ=pB4�TC�����A�,�}7J���P��i5������פ�dg�Q�l�w���:����r<�l���Zm}yl��[��D��n)U����Z�6�����ȣ�ъ�KTe;�e���
�H$��-!~{��9�l�Di�+����Tͳ�n��"�G,
�F�cN&MZ�6��'�F����U�u�������d�}R�_Zt��_~lJ�C�k�Y���wm�uR(��D/��j	ɏsZpr�� �$|'�w�QF_�o�;������>7�Y���V�ƭ��)�1�]v���iP���b{!Pr���`����{<lash��sSk�S#P�O��yOc�<�:P���f��ɀ�@��ҏ����n<J�U�e�jފ_��H��;5�J�_���O߿{{SM�����\���^g4�$5A���t��D�#d�*rD��&�����4�Gե%B�/w)�����(�@�����_Xk�s��2�|e���S�F���u�ݘ�z.�x��Fx	lPH�6ȧ�'��9>�L΍�f�a4�f馸)�ʜ�Ө�s�DHa���F��t����d����#��U�{MA���rk�j���r���JfIQ0�z�������D,n��C|��4�1I��n5�#��"�!�s%����D~ZcH�:ppHG>�g�;�-<L]�y�z��L~��e�	�f�'�Տ��9�zQ��KIv���Ao����wK,M�����]e��غ<��k�H�&��hL�3��)�0��dfE��a�}�,����۾��ɖ�s�3����V�м�( ��?]䕁S���[�̜m��I��m]̥�^�b���z���ك���V�S^>7�+W{�?�ʞj�ꅨjs͏nX#BTa3�ďXgΠ�&��G����	�L⿭���'Dv���,��-�ޒ�z7ǞF���������Y��%�v�,����o�=W8�Ǽ����E�6�{� �."�x!z=@�1\���9�J�}(�A;bG��ׇ	~�Z�e���n�*7�GQ�yUh@߈UɅ���*���P�j���n�C����x����V�3�\���"�B�4ai.�g�	�&����1�׽rH;zK\B
���rĠ�M�Ᏻ��;ʄ����?R{{z�����&w�"Q�=Wjxf���(WB��V{�
�1��Ǭ1,_
%�=̂��k���	���Q��ÊR+��]PN$���p�P7���x��l>Y�`�f���,��G/x)�9_���&T��5;�f�s�Qo@!{���֏��w
)���T$�(YU4��$~Yٌ��z�(qc,�L���"o�e扨�,Ep:+G)n����:e����<c��fQ�\goo�)���/�Q��4oO��oymd�+������IM�QD̎'�\b�y.�[ݸl㉎���os�e��up�[��sHP\�(b�ls��>�~d�4�.��ߚK����Tς���]#�8踏�`�N�h��wG8F緗O@��e�f�����q�� �����n���4�q��lZ<�'m�m�S��7怕0��rE�8$��Y��|���S�}�O"/f=$��v������Lൺe�Ѽ]�J�V��h?�0���C}��+E��a�v����1-I��R���Fv�������nx�i�z�8r�߱��N��q�V�CH��V{P��LC߭�@��OE?�N��Y���߼y��	���	G���6�pe6,���ƌ���"�P�9�MI/�u��>0A��5�}�3e��/#�W�y�.�ÜSo�!`��l�%~��%��ځ:��������w�_HYz�B��z M��xa�	 0۷m�w�v�Z�{T���=�Ƃ[�_��X؞��ғ�zگ��4�gC�a��9R+}҄�-c�O7�ٝ�Цw
#�X"�R���f��������#��p���	of���lߒ=��E� ^_�y�6�_&4���n�l6ky��0���˃��(��bo=7]/�-�PB�
c5��)Ĭr�.=MVR;�&��J�Fw��m�$8o-�@7���� �����[��<:�*���L��~~Z�u�)��9 �x;G��4�[�]�/f-wÉg�~mL�,�d�Yu��תK����$�QX�܏�ua��yO���V���uZ�=38�%�g��{�f��P�wm�кN��e��k]Y�_l�����ZL'��7G(n��f[�'��ɠ���Z��c�����a(�-�A)�$�!Ы3sJ�W��7_�l�$�NѠ	�s���nqG���:�9���d��y;��R���sc0,�kj��l��m�4���p�P�eܟ�(5u)w�*�z��H"=z�u6��1,j�fx ��pc��OvJf����j�=M��2�b���e�S�N+ͯͪ"��}�Q�-�3�D�xjѧ����7)5��=��p��;�}��r����W:O2p�kl�E�<���r�F�	�ɗ�4�7��<���,��j����]�/�O|/��z�K�B���iv���uXQ�,�:8���T�%(�	�@�m�Փ����r,W�����(�}��{3ئ��_V����ě�Sro$�y��W6v��Ӵ ����|���U�S�.�/�@u���ag]{��f��O��m�(lNo�#pp�e*���
��;4<�q^��v]�D�$"�#��J΁�TUÔ~�e�H�	�Bќ"�	�ߵ:�H���g����<�?��y>o�/m�?�"�����KDj*��$8���0�נz�,���a���̀�ߟ�����,xg����<E@�I:�f>���-vr,�v�[��<j\jX�`�hؖ%o��{M��M&�-����8.rZ:2ҹ��p�N�c�JVMU���U<!P�vS�7>Q��H��Fߝi#%މ��Tb���{7���
F�.]1�5��pX�|�w��\��&s��V��&��Hkb�^�}���eM��]���s��q�۪�8:E�Uʰ�75���;��B���Z �.�(FJ�}����z���P4�r���9�g��������2�nt�*g9�bx��Z%�UTQx\�4�4~��;8���M�os�����?fxi��n�@"���/���`M�_�7B��鍬Z.�!�v�<CĹ3z�S��x�च��i�˕��+a?��ż8x�F���Ư����dy2M�|PS����X��W.1��nc�ki�&	��4ZX�)t$+�uc�	�� ����c8���49ş��h�e��D?,��4}�"'�xh��:w	畳�	��Q�#o�����5�'#!(Z�\Gǌ���} Q�%f@�џ�U�9�;Em�lT� å>��]Ϛ5�k+�����ɷhP�F��,����y�fj���+w�_�>�bm���hZ�C�h�#��r�Kغ~-|(��=�Ӳ=�G��a6*����hi��� ���?h�_�O��I��<x� D�Y0�`���0P�d�O���|�w;
�J�g�(�G�����5uѨ
*�:�
�d���0|��TQ9��:w!OQ�Cʌ��f��N&Q74]�$�9�w&i��ES��-a��=���&C�'�B�z���V��	N�%ѕ3���.e*
�3?�6�P�y�sğ�y�� ��R����Q#d	mh|,��\��-	�9ax9/���x���9��=�6Qk���1*u.Li#!�a�	���q~� �Ϩ;�s:����x5�� m�Ⱦϧl���vq��P2�xx��%N�k��|�\�d���S	��h8�m��B�1ٯ' n���"��y�0j�q�m+�*;|{��ˤ4�����*�C��A�r;D���ei����@6�,"��A�d��c�`��3��j���v�	��5�F2b	jM���/��&L�f|�W�vA�md{HR�g�^�qf|g�07�j]�x��XB	=��
Oѫ�9f�l�����RsQ�;�m��`��O(Uyg����ѷ�p��']߶9q�z���3I1��3��x�"d#I�q1�P�gO��}��&j�w���?T��8��pE����n�Fu�~��tgk�#���YM��}_
�R��:��7n����U6T``(�,��+�<#�D��Hr����&P�f����j%�"q���C�]�huX���n���$7����(�>)\��k9F���	c$ٻq>fa�n5�@���aK�|X�I��b��ӣĽى�����6	*X+o�ب뼮t�I�[`��<�*o�3[�Y����ߞ��5噏���zm���;ȸ^�c!�Ɩ�@��vXX�E�w�#��'A��Z�����II|/0�l��27�zZ{���Dǂc-��	H�>� ���ш�^F���> �e]�P �&+b1%X��2 b�ζ�1�Y�Qm��=w��kшU�`��$	<��Y��֒=��z� ����L3tW���6���Ы6�<����bg�X�'�2�~�0l\|�rU��;}Eta��]�őy��o��Ս3����~���d���� U�~t7�E�D��:��*E�j��W�^y��o�����\$��>Q-�+n�v%�*�A= ��ù���R���0�������-;@'���s�����{k���!���v����,YH�8�t�(�x�]���֔{�c8���KW���L���5�;PR:vYgx[��Y��qM���Gkak瑱t����{��~�5#n�ge:2&i`�۠R�kT�\žY�g�9�K��KW*e<��-�-�z��ۖ��+��N�����.K,'?��g����	'A��=���!_6)���k�>>��U��"�sby�% 7�uUv�m�$�z@wF�L��q[*�COm�Ac����{�P�pt�1�Z+�bu'��:�[ݦذ�Y}�͝���/�{��݃R�w��?j��.NN�k��gQ�����Vz!��}t~���ؤ�Y�c;�ZS��d���D@JvH}��9N�� f4���;����O�.u�˽U#��h̠0��z��d�pz��hV���� 8�!
[��Q6�l�u��Гz�D&h�&pѓ�t^}��m~NX�y� ����+6v,]8Iъ�¿c����"��tW���(t�;ȍ���&�����[��O$́�V��F�guQ�14��<>�����B(N��tT�A��(��b��1r3gj)�''f�̭��v, �*�ҏ:�2��b�P-`k���{5��=�r�^JDKV��{��L'�l��H��r''c��fZ0�6��F	�g8��������{����Z�XM�����]k"���#�lN��}�V@�U�A�xJ%��n6J�Y0����4P�D�&~�ǯDʃ���g�^j�D�Xם�ؾV�~c�ޠ;˚׫���F����E�N����2v��F����c�����Q���_�w���:߱����	��l?�v�����H�v&j�&4o���~PX��Ȃ���?��n��s�&���g�i��}cHmy,��I�gQ�
&��^������zu熇�}�T�B����G^�j-��[�c^�x#k����E�J��Iw��(��#��3��\���̾�^)_I�Yd_OQʏy}Y��X��AO�P���Ip{M���Q���$1���dtN\��!'�Ӻ~Z����/L�T0�|�i&�"��1\���)o���=�·2뚺M��R�~O2�hil��;7d̿��1{j�-������8�H[�bs#V���d��CZx�՛"���q�jc��	�6:/2�ㄢ�"���t$1��B�	���B��2�=��nos�G�wib$���\��;�����b�D��u;��H��A��)����;!�E���"K����ZB�-`ʊ9,iz�g���lTB���bi~. ��AI�,y��eR��HX�ᝑz2���jUgimy�������P~hm�K�]YaL�w�+��2�ѡ�K7;a�!�NQ�Ez�:T�"R9���k]�Z�RƳ�:�AP��P�vL�΋ԕ�;!WU>���If�,	�٨� пt�e��_,�̥���|��<����o��<��+(I���"-��esf�2�Bg�vb/Qs;c�M�tY�I��6��gK�'4�J�[^���������ބ/-�Y�b����f�z\����o~(��EaG�-���9b�o0E`4��z7�uLg����f�
�؝�؝^k<qD�Vcmx޾1J�-�u4#�;��u�h5�%dB���ݼ� J2�z_lħ=G�C�ޠD�双zB��l��Vg��W�����@YQ�s����ƒ���J�uiV���T-�w=,�zD#��5�֟�_�ݐ���B� N����՜���tQ�ڋ�,I��
=��"��n� ͟���쐭�ϔ�oKT?d�&�Vsi�N^'!e<]؆z0��0=E���j��w@�)s)��B~*�b�����v�	D%땭$�R��(H�ɾ���V_QxM�@�`Ft�d�i�B�J'(�kM����0>R�=�6ShK��TNVYk:��l��ʝ����}7�%BR��_�&�au��W�ʘ	�(���9&H�ףV�Q��m׸�U`����_��	�����U ��TQ`�*���V�/� ̸�!1�g�d��!p�(��f�i�b)_����V=s�}�irT����t����6du2QNaʻfěL4$ꂊ�P�ѡ�W�bT�R�6~)���b��t��N��V����H�T�g��Y�
�:��P�:U�5.�A�z�����Y���]-�B�Rp!�O���қ�4�����g/�2c#w�sA-�:]X]sJ�涄_����Oܺ�E"l�G=�U,��,�r��N��
��y�7�>�n5�������.)/��M����a$��$�yt���w&:�mYS��٣b�\1��Ey�3,t��$2��n&�I��Ԁ�V�;[`}�A��C�����(K��v����ҊA���}L�~&�V��p��Z� �Em���{g�����O�"�C��;uyY�ޗ�GNUv�H�92��pӺ����mE��0���%g��`n��ǿl�$����z�7@�� ��b���X+ͩUi�k#�S��ד������}�F��F���;<���.�'�D�f��g�8֫��	a�VLz�0�T�Ӻ�r"�;�?W2�=My��<��W!p�5/0�e�z*��ˀ;��W��*��Q� ����)�25.�ziq0���Rj)+�o(�#��DV��`tz�cU(��l ���'�f*4댞�g�N$=� ߽͇�h=���s]�oٴ�yJ��m{�S��ʶ�~2�}���'ȫ�HdFҌ�[C[g5�V��"���|�A�]�+F�6�`�h��.P>��R�:9����f:�y�j��{z8�\���=i\1 e�1Ö�����R��e������,=�>]4�"ew\ߛi*��3���Oѳm��9�TMZ�i�̰�s�a���i)�6�4s���>�1+� ��b
P���.	� 47�blݘ�Ui4�͖3�DW"ѭ]�nPF�H�+�*UX��x(u��;�췘&g��frG)b�dOcp���4pP�.�PbZ{����ȭ�)�b�
&Pj��2����L@�� �璘�K �
CL�`�㴬�|��ʦ��bW����� ���(t6AX���a�;�Tp����"���m�꧰���5X�B~t[�L�hB����j�˶23��O��cͬj���2a�=$�W([�M�Db�eO��aH�O���$��qJ.]��
O(
����bG�{�[Q.P�4���"V]i#� ���_��A�p��5qUN�N6r����L��'�4yJ/y��0��"�E�$u��z�:��_f���%~dEy�Wg�'�gb]�`�����
���WV�7%*�'>�.�A$.u��k�s��G��!�?i��UZ�+�	�{q$�Ι&�"}?��CC��G��-CBWX�P+�l�1�-B�0MyU� ]m���f��6�=�z�	���DӾ}�G
F��j�S�FR_`(�G!vs։eIņ���ۢ���Y�T���em�q+[��
�vCE瞽���P�N��g�c��BZt�_C�KKp;I}.���9�)��EP{�Ϲ���d��,����f:yޱ��iŬ���u6U/씀d����}�n��O���o���H�Ca(ގ�O���yp H�ߥ��4�ű��J{�7I���V�Ψ������E�i���]��,������j���2�������>� ����ģ&�ay���I�O��������5�r�yyT�����L@��TfS��>f,\ޢMc�Qe�r�n�|WY���t7t8\\8�lf�	jT�J��4�X���t��%֩[Š��W������f�,@ui��_��*d�a���7�ȧ�[:V�h��K��<��ޢ`m5I����z�h��/�M���|a}�R�����}Я��<k�Ȋ���PFe�*>S����Q��&�M`[C�q���_�_ @�gG�,�0"���ߡ��Gq@4�>�ae�[�=J��T�I3�9R���������j�HoQC(�q-�d;�Һy��fi�9�j6�}��4dAG��O��e��M��[K��� 1�蔍6�5�7
 e^��CB2�h
3����Qh��S�;�^KXֶv�:p:ɐ���W����%�R�m��b�S�14:�=9�˴C9V3*� ��th �f>Ιl��]^<ߏP�L�����iֵF%.�`��-���;�����i�&*M��k�ut�M�{F3�ezq�(Q4DVa���ş-���9�5m�Ԯ	ǉ��R���G�C��!rk(y�'�d4'��3�:vdǉv��o#��� '<��7'o ]*�!C�qg�j+�-��ϛf���ޣ�/�#����5�V��(�" N[%�P���YNG�#E�ι:[�=�ەƲz'��@N7�}ޣ�YS.�.�W�T������]�������>����>�B͉n�U<�n�d߯ݒ�q� ���.gF��Y��]Q���}��Gm]q@�n~�sy(��K���n�w�l�涸YX�"�E`-�c(��³f?wR/43"0�q�
�TH�-����\�� ����LEG��*�����$9:^��ݎ|##�F�;\���&��1(-�@�)2R�$h�nlKc �%���dL�`랾��(1��I��v7�����l?x:�_�/�k7�~곓���,
w*շ6/'j?�r���b��Gqק&�;����opbEb�8+�w�.T�=8EJjq�A�z�;Jg��" ͒g� |��P�T:,y�4S
��� ٳK��ֽUӎ���{ލ
o��G栏;x��R���]'S̱���5O��7�B[/�K�0�Oy��J,�	`����Ӂ� ��{Q�_}w��pϴ�`����`������Hc+T����S���Sk� ט#;�������DX@{�V�+Ab�"-�Em�jkb��}�n��1�\��C;�u�#����g|Y�5��`��������8��Mv�D��'���c�H��9���H *?�a�cJ�����e@|�)�ɨ�t���1����U{i�ch�K��	�դx�4{T�%�����yV��r�t��+�_a�s��3dՖ
��M>}����-�H�ݔ�87{���*RW��MT�-���U�74�<`2�3*$ݳ�;���씷d��%�t%�:�BNc����V�[���-�c�����(B�K�]"������c�
Sog�<�2ī]/r��ⶁݮ����#	K���?y
�٤�- '�H_>��7Qͼ�'q/2癆�qB��S[:j��E������(������u^�d  UB'n��������:ly�~�4K9�Y*�,@e���'|r�9����7��fZ�:L==Gt�#%Qmc�(�'��ܼ��訨>�<*�VJ�D��kV��2�;�;Fù��4fn������g~�6�]d	��d܉:�������������{n���e�{�P��m�D��1r5}%9��#gB�JY�	X�>�(�(+5M��R���� N����!�UG1�X������[��d��/��1Q���.��0��a�3l?�]�T�4�O�u}K�����I阮kCY��x������x�H��R�v��ý�~�S�ť84f�+PT9�	\d�A~>f"��?֓�c�� h���#���UKј���&�� �h��
��qJ�H�7Q@^V�lLtwJ�9�L�b ��Іw6�o�k��Q�s1X�b_�.�L�� �N�_I�e����1�`c�M��<?`����	��I��É8LEd�ZT���K�0(o&�%���c���2�2��`���}�r4��}_��v-��J�OF2i�l���`	��]�)�%o��1>jK��Sy��F�?j�����m�,U���;|���BDa�h��z%�E*��)Co���"8��t���X?jAJK&��RX�6��[��M XL��aۦs����i�&)U��D|�B4�d�I�xF������}%�.s�Xr� *�/o��m�MLe���F賗�D�����pL��o�+rc���g�?�N3�V�K8��{��܀q%��]�fu�j@`��uY��k#cM��Z�M�:��<��,E��� �æ�V�b��6N���M�S֏a�T��ؓ`���ZEO����ã����� ���L���V�¢���܉0�m(q<�kr�*��ϒ��p�(<���u�6}ӽ� Xpk�Γtoh����F��hh�0���)K��b���ra �:թ8�˲ԴDM���H�dM�a�u�H���� ��xL�`ߍ�9	=��
�g��SC)$����c���%���L��h-�"�Zf�`��a�r�]8�ߩf�2��	���"j:����L��hPt:�A�"���!��Ј�x�.�.��wU�WA����œ��
Z��7{� B�eA �O>S@\M� ���`[��|�={����<�w��� m��.Q8i~�*�3�����b6�
�[�˔�%C7�{�V�R�U6��n��L���u�S���M����h��O8Ҽ����^���@��צ���]�z�g����.�2x��	L�T�	i��@�����p;�-��G��z�xg���8�L`����,�#������>M��A�[2��jK��
tY5��A���(tC`�J7	d-�?qy���e�������)B�[C��Tްm�LV�?H ,d�ه�E��:�5U�ݘ�
��[8�iT�+��uA�~�.� n8����h��O�G��ė�hnTG#g��3�Ϊ�>�I�*��P(����J60��@�m�(���P���l�]���J5H��e�W�ӹ���.f�i�
V�%H^�J2�����NvB�7������-���ә�y_�����NA�z� |��ث��W�n�N�s��!�$g��g`s��<��>h������
�s9󒪝S�j�� iC�Z���o��x������r�蟪�+KQO�!ڎ��  - .�v��\be��O�?q�܁���>w��cص�8�^���?T�O����a�/��Tc��~�J��d�[��Z˼jdA�C!���?t�:��BȺ[�R�ut��O��o�К���8�EM{z��z������/��S���<���F�a֨h�[��JFN�I�,�d����)Y!֥����NYv�B&���}��b�E"��?����:�Bz�
�R���?���ۡ!|��?3b�Jzf�d�;:�6Gyq_IpCm�p��&Ʋ��P��$J�Ҹ?I�I�9p����Ɏ�q�o[���>tV��{ [� ��M��X�"�c4�8ґ���(���XW�Aί62U�e��;�FD���Q���a����Ai���5m����M�nA�����O�o;�����,�� ��ܮ��|���-F-�`�'���<*X��w�x�W�ZR��������[i��k�r��L�'y��Q���=��h|$����o3��/TRI��v�?��n��D�^{4�׹Gm���,���G��Aq��g�HSA���T��/�7։�P@3x���6��7�fFjC�8���_�1��D�{]9?�2<0^���N��I%�M�����&Ƕ-f���������3�p�%�9��!��V�#���E6��v�z��>�(��w��+���ly�u��/��ܾ�9 �k�e����cH�Q?U�H����P�/h�b��u6�J�l�$�1��_,rA��D)5�0��d]zi���
Ո��?���r��֯�'�5 u�����*�H�����
X<8Q�����9������=�ppnӶn��0(�W�6<�+K���~�+>�Tи��r�z�{l��_�N��Z��)0�^���T���4!AE3,�g}y���ޝ$��6X���T��h����{%��y\��N�҈g�K�ڴ��j/��-��qiIFCc�e��@����C&�J��Ϯv���W����ζ�xP˼�����VI��R#�lR�G���Okjqhؗ{\���TՏ�M��,#�9���a[C�*{�"��RjG2�WW��N�<�-����*%�Q\$�.Z�+Gy�86�F������p?����rUE��G(���}���=�X6�9��`�����V���"��@��p�$���Um����gw�T g �k�<Z�̹b{�'��N�������V4�ɚ�w�yaLz|�q�]�ݴs� 1 6!����F,�d9ϭ�%`���}�!R�$ah41X0�$���E������H�7�TP�����qgB����P�	kDLry���E���W��B��8�0�g�vj��~����T}¼|�T΅O���WӞ��ǋ��8"�����s~Ţ�`Qo`	������N|��Mx#ZBۨD0�|�՛R�t4K��~����BK辟ё���,���Z��^�K����G�.��������
�tM�I���O�P�|�*��������fk�������y��n�6%g �&$Š���z����A4�9jǯ�.�,!�ɦ�$є��Q�{�d��Ӟ�_��ڶ.��*�(�(���H��(�K)Y�/�".���	{�(�f��oy!T3����F}A��2�T�聰�cpU��^�b�M�T�ؘ�s������.�\��[��%����{W��	�b�봆��V��1i���OF��-JB\S�6����D��8�x���f��� �i�Cl�S�apͷW������_�� $+X=O��&8-T�`���R��jS�ڕ*�鏘�x�")lY�՟'�؆�g�f���7˷ҝ�#Z^Z�£�&�L��l5�i(L`��_�Uҿ6�](>�_`�T���u4�1%�͙
��k�W}>�eR������B> �A�Op�&9�������'xO*ɂ���H����#���eE�G�*R�"��˻Ǭ�5���R��
�X��5XcI�j���5`�4ow�#Ĥ7K���.��B��U��I�Z�](l'y*�6���p�$�G�po4�cQ8n��w��*�;������Iy;���X����C���|7�k�t[`P�����MK S�!�VLZ� �ꙬR	�����<s����c8�@j�C�#�h��@$���1�YzZ�v��#X�A$W'�(D�a`�~+�_�<���R��^O���ȥ�Y����]����VX�`�e����"hT��(Fs8LPa��x��]���܉�[<�*Mv`Z�Cv'�}�rj�:�P��0Tȶn�p��X����G>��ڼr��Y�)�ۻ\�w V�OY^d�'�}C@�A�gS���W�r�u���RL�6x�.4^}�r�cT1�8l8�_=;���A�/"���e(v��i�>&�/�.�~Y��2#�}������ݝ�0�~�L������P���D`�e{ig{�@W8u
G&�9�& �%��f1$�ޝk�㷀�lȧ�D���d�<*�l�`�q���b��2/v!�1�,��}�/F���Ԯ�\�˝��a��p�_��f�̬rG�u�:+��F5��{�����O5����'���E�#�(��y�"� &:P���:V�A2Q-�?��>{@D؁�}~��A�L� ��X0=�ҝl��S���/m�v^��wt2�k��{/Hr[��#��=!IZ���F�b{i��C׀���b6pes��hh�� e��Αϒ����6|���ɢ9��O�/����bs�I�������Z��t]�Ò_�~����&�3:V�G]�dB��#�.���H�ͣ'�*���Ё��oY��̈́���Xs��~.��p��p�,�/�&Ϯ�׮�բ��YP[��2��
7dmR7Fj��H�%���l��0`�%��b�!�Uy���5?Ed�w2����?�����;�o���5\7�N����6�ջE/-D��6��]g$}-���;�zi=Diy��f���A��q���2����x��g�}��_f���0F�y���Ib=����䈾���H��A�����T���/B.���VS���SH
p�{��#:lzH:�����G Wo���",
�#d�u�Yj�7'?c�_��ZU��yǬ��	�MyNLdT���z�a�c6 �E
�3�^�2��d��0ht�eBS�i��g��ͪ�x!�ÀZ��wru�4�J��h��NUI�D���9������������2�xpfAz������I�>b�IkTm���� =��찲ǸX!��y�]7��ܽ�o�Q��_�3!�U~A�+���"ޥ�{����q��u�; �y���#-� >w�E��jw��m��}- 4�6+�CZ���8�������a�:t��3��?2Q��C�H�H��� :O��B�ǎqȖ��]�䎿N���� ����Fd��Bn��p�r��	��b��4���W�w:�g�R��O� Έtkf����G�N��\f^��uǪL	3�r���`�%
�����ֆ�~6j��8z������6o>V8�r�	㙪Ը�նg��#�ƕ�%�o��=����F�Ñ(��Ȃ똀X���,L^$�E֭}�˩�-���/��{�0�%�d�����`UIYA`�<C�b#0H�fIaT��O�u��� �)̉ށ��~\ȯQ�P������E������g���s|��Z��D��84�?�l���F<�
oD��sR!]�R��6aiCeZ9&� sY�5�tZ�(0TK���[.u����ȑ�	��\�|�*;Ҏ7C�uVj�a����fq������bhm��e�lt��R�'�Ӏ�5�e"U�ɇ	������j��7ge�
ɒ�A��ᙛ_�b2�p�㶵9�b�[��{."��FZ�=|��r��֗4m�k1<�T+u�^��l����aW�ѧt+�������$aD־��:��I����n�m'�YQ�|����(?IZ�
&Q^VU�ʤ�QȷIVi��KtZ�k���o�� r�n��eݰn{���w�e�cgzj?E,�:���Q�%N��z`�#�H��Q�=b!*$�#h �ר����X�:�����	�W���;��һq(�"!�ν�߮I��� �Wy��yZ���=��p�A��~��F ��|i��շ�q�l�K��P��jP�3��n��+ݍ<_S�~�y���=��m��[͟md�g�-0 C6gʭ�J������m�(��W'�d����R�ZԀ}rA6St���0��Ej�z/F�g�`u��Q@��J"yk&j�Uf�+��mC���
�`��Em��>��
U�6�T�=4����@=�o}Nbk�
pgd2a�k�&�(�Ꙑ�1ؕ�&UZ|�?��U�T�q)ˠ��$�&ig;����6��C�(�e?Ю�	20[/l�`Zl��\�0-4idv�v�i���q��>�y���B2�����#���Lnj�x��G����g"S)�����'Kt	�ל�5� P�Bb�G:�u��,�!�I��ӡ=�[ ����<lԐȸwɬ�~t^�l��t�t��)®`��1�@��kn�x��p����j�:*7�\�S�A�}�#kaCP��8�L�x��������(�gz����a��Y{��.�v�Wz�j{��p���4���̓�}� 
�;�*��<�� ���<��a�����w�[��צ��yz�0��+ī�k�&� ��J��.����ȏk"���BQ`������W�'����z8O%�R�i`��o�Dռz �4��������v�m2J���5L�<��������
����$Źң%6�7@#��\4��m6M��l���a�2�f3�Y�1i����a�{�}X3�L��:���p�,�B��OXx�(;��>��q\4ԅ��`u{�ǜ֫Ƭ��W�"�j���hߐX����sz
Ee��v�������fȸ,(`��	��.8'�MSb���Q�M�`}P��'���P{�O�J��Hd��(������:0���#_����$¼ܞ1���l�6@|D�W%��f����-���f��3p�h}�*J#?p~�m�[Yc���� �2�Ԭځ�b�a�l����ɷ��zt��S@A�#<q�7Cv�^L��u5���Hr '��!Pΐ4g�c���{g��NȡW�!WCH����4������-qH-���j��9i��~ᑇԝ=o�後P#v��*�<V��`����D(-�_��bZ��RU���]+
S��@�}��ٸ�a�ts�"�}�]����	R\���R>���r�>�Vu�Ks�:4�H��S8�����_�H�һx�W���~%C���rfś䶍z-ׄN�|)g����i#�g���E�H�2Sw�_���$�̭y��H�!t]r#xl`>��U8�Hs|E�ÍVv���W+���*��F O'0hbO�eQ�Δ'��{�.�DU�1�>��ϣ�c�9-A���a!'�ٹH��.��w�]K�'Y��9J{�ـ��͡���J���F��9��K)@�qb� ��;�@<t�GE�!�
"*��c�O�����,}o�ez���I�T��`aT���P�4;y#u R����?�� b�g��v{ 	��(>Zmi>F,C��Ad_$;kK��y*�[�3��SQ�}nִ��@�sp�?;�THLKo	ݴ�j2om��z�ch՚��y~�6�K��^����/���&޾I�`
<+��z���#i�^sj�cS���2H.uL�V��:ʕ��7(��'�{�	�-�F[g�G��hڛ��?�ɚ���r�0��x�(�~�:	�\;4�fp�\N�ec�E��U2Jo�F}�i�����t�MIc��X��B�u���7�
��737�ևw��/�*҄���:�e�>���$��m�^����G#��8��7�\�^0sG��Wٗ";���<?�&Π�&r�F�<���Zb����Ve���_f]���G/m�>T���e!����x�RZ����i�%^;���Z}Y\�@N�A[�U����\�7��Sy��	�S�D�"PC�ڕ��-!�ێ�W�a(���G�.���o���>�V�K ��������%��wK�}ZƦ{}8�3P�2���v؃=�L��]�Z���bd+�Ce��ֈ͝���R�'C)K[;����x�z=��p�\��0<i�| �q�L�$=l�Z�u�NKG&R#Y�W�z�/�6��Zժ@A��U��Ff�gt{]�R��̍����I	jΚ�7LzF"h��������Z�ME��#:���i-L0?@6�Fyn�d��J&��^�|�]ъ��,1�ٳ�9s�y\�� SR�Z|�U���m1�e1��'�Uaٮw�i�q��l���z׆���9y 2s�E��6T������5��J���3��(��(��j��;������L�2"���/x&�~�P:��<����1����@"NEh��J��/�J%�	��k'g"w�ú���!��6��h���$�į��)Q���,z��bE�!0|?����!u��:�6�Q�XB�o�3��Yo[�5�3�E���l+��GS��lZ EF��p��^HM�{(�n�"��'�
Q�WtSl�OU��脭x��p�a�x�I�{C���3k��.�� 9���gsA�,�j�~jF|�IeNM�\�[|](H�'�ـX��tZLO�����6KH^�6Ԩ�B��'�!��������]�iх5�a<J|���H�A�9�K'���ݥ� >V7���<p����'�^��)V�e<��^�B���'���� �W�Z�axG�G~��"����lu*Aj�N�qad���oR���YTx��\�cϔ���*��]��p�:Y�fI���T�}�c��`��,�����lC!2�i�1�D���+�*���Q/i�ڵ{������P��"����d��k-�}]h��uē����l@��0ĸ��#�fw#��G2�A�9YA�נ"�Cy��wWH�@���cY����|�PO�X���YTm1����_�s���mܻ��_���
��r�N�*�Pɪ�\�g�v��-���4+	$�Rf� �W.�\vAe]V���z+���ʹ�(����{�=4&����L�t����?���=������#A�٤���+j��`x!�����L�gah(��+��z���LB����b�r#A�'��8P��|�ɮ�Yb="i�o�^�i�&"� \���;�})!�Uq��-�
����QM�_��Pn���>v�pT���H���.[�B��	S.)�*���Ye��yӈ+���*��Y���}`O����$:d4���w�݂��Am�֡�:�i4w���^Ӏ_���m��wN�r���JO�ˈ3ӥ5P�:���u`5��<^���,�lv����ՙ�,kN�0@��|P)��s�G�<5�bINP`��l;t�$9��ٮ�_�r��=c�Ά�8y��h��X�1�yc�)�-I���c�>��7y\�t�5�F-���Oe,V�U�;&8��@�0j�m���z�5Z�l%	�ϗ��S]���wO([��IRѕQ۟X[܉�TV�u{�����o�K|b�f���J0_�3=��ka��J&�K^��%4��SN�U%�VC����4]�S
VfC�ޒ3?�D���*`�oz��kK�a�����������,�,+���%R�F1vA��5*��f�L?�����o_� ,<���k�@&!�*
�VAv-xN&������1��:)&�k���e73�����䜽a]�R��n�D�+��,l:�m����Ά}>@j�d����~jw�;�0�Js�\a��LL��-ӛxܳ���|fpi�y�V�9=��i�c35� ��K�8�%8u�h��Iѫ0��h�r:�:,u���d3�5Q!��vu2Z����4,��Xrt�/���W6��<�e�?&L�.�����(dl��/�e]Ѫ�Vtk��?w��ħ�v�o�����%�7͋���XE�6�[�?g�.���q������1T�.��4�{<Î8����qH_ʔ��]�u��d��%�V�_ϸ��<��Mܮ��\>�~R�ւj���
ё3?����=z<B��m�[mO�"n1�z��F^�(����=Hz�+\��/8�n���<���,��ާ��ظp��%gY?��Y�i%�&����˞Vw:ͻ_�7f"�"X��8�χ߹�_�=��/���S����;\�Xp��9���*G8-h��aP���d�C	����>D��s3Dd1s��p�1w$�˙��~}p:��A���:���`R^�:�j�b�)L>{oS�X� u0;3^��5z���^xWݳ�ǗK�á����̄"]M�:�����
�(�Gm��������c�f����`�$�T{KY"��Z�㡒�o]M0��<�&��D;t�&�����գʜP��d��)���}6%����_ԃ�a0;|]{ڿ�h4	�l0#��z�$b��o���H\�m���l�oiOsch+_vzűO����`Gw� �ض�=xY�`*��B�vz���Z���9����ٳ&��_���6geF��r�:��*�M���ƅo%(1}qSS-����1�l���^��7ZqJY��y�_�#9���#;{�½���-�)rE�w�S�=ܜ��o1:?+�Lr��J�n�ϙ�s�1�����>ˣ�@�WELe짳Л��ҵ�#f��W�/�E�?�%�@����Z?v^ d��fk��N��r����-�P��!��R��@�rs����^��@n�����0d��3�1
L��)��n:�,V}��8��E�s�"\ǆ
iy���f7r9��ɵo���GM,�}s����QȣA�R����Y��-POG�׻J|=Gؒ< ��o�?~�D��2Q�D�=�?��ܾ���~cO�7L��>-����N@�vb�,C�J�ƶP[���a�Ά��+ ��`Xf R���
�M�T�RNWI�8@w]��|�erh@Y[<g�9����w��"l�<��Һ��p��O����d~[?�<�.v�^7�(7[���A�J�	r�jY��|GuØ��ɠ� �7��8�#T�MB;�P+4�ji,w�.�d�hô8�Y�'??y�����B��S��)�tS��,ʪJj���r�K�G0K�.��ٖ�ĥC��g���l7�ڲ��V�H>x�|ק8�!J�����pe��V�·t�V���{�E�G�}j�9�RA3�����tn2���l���Q��}��>2n�X6�����N��K��*nۖFg�;�tNè6��P��q�A�'�/o��
Dq��'��G9t�2�S�w�j���w���QWd�Fd0|{e��c��IKb�����i:*uZ�>[�h~`ˡ]��2bܾ�n�H'̕d����qa*�n�շ����<s����v���eb�¼��	��"|P��!��br*��Rul��}�b%�KV�MPiJ�CЈg�x���g����=��8��@C��-<���j�	�ɢ�Q�*V�t���aWv��� ���
�;;Z<�p"�n���7�I�|�����"Rs�@4Ȃ��:���IK� RHNDY2�`�W�H��i�� �c�������>/�R(��(�x�����: ��F-%�$�MZ�r�[�u���R���z��X쮗���nat�/t��'�ŭH��d������պ��a�mfPᐖ�>=�O��z`�jV��sF)�-5�.�y�<h� ��"	K�%
��*�+$Kͱq�
���n��j��}��g,�@5�K�����@=��/ ��K!<t��`~���^W�Tm�jǹ5�u��y�2�r�D����,m� ~g �yb:��s��8��;y�IzK>K�Ze�6�r��b��YEV�����eG@�@ʭ]E�FU�Ye@���)6\b�u�m{��z��3ʓ��.����I���'�J�7<R!�"
����Y���D��JѦ��*�w1��J�|?n�SfU�|�|4)��������a�ѣX��6 �M���g��Ũ�x�і/z�lv�NVO �o�+�
��3m�U�w�gMs��h�
k�$�}��>���>�³�-��JڮF���zX�d�(G��V�@�@ĉSnj��xK|s��M�MX��ȵI�x�\��UG�_-2*�^��L����ل�o��C�w5S��Qm�6�T0�ea
���(�I������u<��M�l�e#<�0��#��?cU�;v#IK/�I����
��#0�{`�5ʳ�0��؉�юKE�/�$�-�5��&@{���}��|�}@����_����%�rc��\�eke<����,�����Q!��
��.�uչwF������Ў��+�f��)��m�BRj��t��%�e�7#�{L2�ߞ]`:aAכֿ3���%��K��+ꛄ�L��BU�'��m	�g3>�Q�I-zjh�Hh� �A�e�[�U�`��K��jT�
���=fZ���Ϳw����������~��� �Y��'ڿt�=�
	/A��h� �;JϪ�F���+�,yO6:�X�D	���hӋ��ļ
���2��+3 �(\/���@T�[���g0L+�i�2�`JvkZ'�Syv�M�nb	�@�}�j^��%��#g��l54f�M �F.}*|*_�[���:uQK^T��o��&�;ҧ7k�ť���]׺��3���$�>l�H���K��;g�ְ�)ioL�O�Z�e"�}��k}�����7��,"�*2�:��b�4�����'�r����k�����c����Hy}�F�4;��C���Wl���||%��{!�sL�
ޱ�����(��Ɵ 2�����ѷ��vj�b{�!G�9O<Ż�Wǝ�P����	<�Q�@M�Qj�I���V�ؑl��tS�M����rP|������
���ڵ�IJ>��g�
��S�֞���Ĳ��9~5ٱ=@����T��\s��O},������0B[��-c�?�?�n�Z�ޜaư�xe�`\G��hv�aΕ��^�$��H���Y+/�!��)�Ô'J�r�|k�A"i�c�k��G�� �*��c����W���j�<��+aztC����
�iY%T��&d�$��F6�@]Y��k��i�y�Xe��	�c�h���#�ѿ��u]�0�;��K���[I��������Վ�y������t`l�/J�Һ�&�q�t�5�Hc!�
�-��̕���1"�s��Z�v&	!D͖��u����4� ��#u� �␤Q�c�a�}Ɨò�1�&k42����%��̾��A;u�k`W9ɹ����7�Njȑ0�Y��B�^�@�� ��琽=�$��H�U7��;������'������_f�����}wO~��;�7ل���C���v�:�35�[��mѣ($�ŽS�a��WY��*�IY��2�A�;�1��QϺx�z����� ) ���7O�j�hh�#��S��4U�嘱Ԅ� b:��f� :�;��ţ�7�^t_׻5iϙЁ�n���=��" �J��ϐ`�8�s�X߉=�Ҳ����vk���L�1���ag�*	Q3jEE��9�(�P���y,C�e���MO+w\��p�����;��4�滵m"d_�?�q�Ē����-��y�3+\Ec�H��C�"+��,$������/�A!��ƴ��x6w8���r^�ũu���{;S�s�6As�@�ϝ��Q�_I��y#~�O�"d�R�:��b�0��
�;�q�d�k���,k�"���@�Q�7W�߫+|�V����tG�����k3O6��W��,{�mq����\�&h��!����źρ&_�F���,��\:�M8���&��Mx�%D.�h:#q����ɋ����Z�oxA�,Āk�g�H6#7��=��8��:w���8�)ר��?z��h�{j�Q�	�C��R�f(�a:L8�릎Y���|��=k=v��� J���� ���{O�t(�P�z�휣NEA���`xr���cv�i\8_��\h�f��h��\�7�\���� :�����Q�p�7͕R���,�@2��p��'��_�g��W+NL�U:�i:W�O!��SAh�i�L#z� ��.��VY��OY����GԗT�>����Q�MĖJ�~(ZLZP	6�aT(��瓕�K��޲�{��K���uγh�Wsu��<Iʛ٨�$�0h�^�:ޞNWTR�?I04�aG|�۸Y1})U�o��=��Ru�o�=�}5#�b.\n���3Ÿ��6�.ШFI�,����d�w�pv��YH{�C��x|d/܋�/Q)qм��������[��Ժ�e��焍"I,��k@���F	e8b����O�)^��eZ�8�+�r���!�SP
G3H"M<�U��	#Cc+�qb[��3Xu��D�<�]��
R�5�BW�M�M�������Dw���)5�x�I#�͛զD�.�����mpC���Y���3vg;�FZ/��u�'P����7L�_��?Y� �S�^�aN'9�)�j�<t��p�����,[%Bp23�%"��I��a^��4���G��%{�Ќz�c�Gb@�`�O�[�D����
�@������PQ���U=I_�����4 :�M�A��m1ThYD1<�����|N�t8Z`����>�+�n�AS�f�"hF�q�r?�(�ر�C��.��}���q��I�gja�t�,y�
�#�G~^^;����O^!�<UZi*�9v���	�ުeM�hHآK.�Vf�M���n��!���J��.���
�Y}m����W�-���ǻ+������j��2��Ɇ^q��>)�ł���2!�B�/$�y���o�R9�sU�F�&�%s8��h�wm��+]͸��T���/0����og=�f�cHR��B��jDt�
�&(��\xa�}x���ibp7�"�O�炔�(~�{n(������'�q�I���r�hT�0�/�ݞ�*�����f�������L^j�ԑ˵��l3�-%`�o4�P��P5�oćq�d&��t�����Ic,K��bDA#ƻ�e�f|}!C 1
ץ������E��^��$kѻ��v���)/ْc��/��RR�n�#O�]�Cğ�~���J��?����o��4�1�FʶJ4��0��t�g� �#q�"��ckXྡྷh�֏k�0����"�v�ߡ{�<�9���'��y��{������j|����߆U�J\����ȇl���~n�g饮�PE䧨�Wޘͅ�Fbu����S:QA%�U���Ϣ�6�5�;�Y$�H-��]Ud��zG?$��.�P<�O��c�����,H�cl�'���az��F�ޢ��>Ն똑���?LJ���-[`�zPYF�j�9�É[�T��(�|wX�J����!E!�-�\-Y�q93��F�R���?a$}C��<�?i��������:#�l�R��MgdTL�d\�t4�xp�nڴ�ǲ��y+�
4�3�{ͻ�?�k�iԉ����(*/��U<�G�^��� 
�Fg���r���O<X^����F�|pL8"���T�W�e�`���V:��n:�9�(�9�vv�1�5s!�v��ݘ�j��w
���T�=��1	�]�3.���V�Q
AQ��t�P���X� wx��#\�gGok�X\�<��%Ipl�APw�}�~�(��˃p�|w=�\&��r����έnb��,��!A������#�3�F���4�O�v}�V������rJ16ގ`g�0��E&Xbl�D]OGe&g@J?yX(l	���E�y�e��=T��*�l����Z�6�>osA�J��cD��1�j���	|�Z�C+�% ]4=_BT�c�P�r~,�t���y�M�=���9S��Ő�4��I�+X��]�� ˏ�@��)�l�CΑe|6��tm�:�-���)�h����|��8	;�$w]MhW���xX*N �k���q2r�d��Z�[�{0ڣ�(q�����o��m���ȴ�c�O���r|Oqg!Ѡ�X\�`j�>:����W�^H3REh�/�"_x�X+7�B�6�#���)KR]��H�=��3�A�P��KLjH�η^��Ό}��ٟ#�զ�]����G�!��I4���P��2�)���R6�Ugn�E��ij��"'$
�7�[[X� <ue�:��
��(V��x� �+�!#� G�p��d�V�-����辉�*��1e��ߜI�c�L?�/��iK�W�e���M{�A�H��eVp���L-E�P��6�]h\a�����n���юد"�h���m7N�`�/����}��). �ܥ��E�`q�A�"2GDܑ�Ɍ3N<���X�@�aP��n%���{�[�%5"VH�ԡF��)�^3�oT�W�ZG^d)ⶆ\4�~�A�d�H���"t��k�\���e��a��Z4^�!^R^�[7���r�!\��7M멥�u��HX���jvVDCoוy$�r�ڐ��$�_a��b�b��0�l����˷�0N��J�x���Ⳅ��v��Ӕ�T�hS�8��� ��M5~<���l~�+�3�� �િ"^�K�p)X=���0�F┼���R�f���J��Vy@�X�.��xj��NL�YPE-f�������#��`��z��k�������{V�B�Bl7�1Z�O/�U���n�� �W�h�Og4���5u2
<�|�Fj1�a(t[+������r�&l�d�2	�f���򁱞f���l��lՎ�Q�U�{�:�&F�E��M�0	d{.�u� ���������[{A�ox&��;�~y���՞'�z���I�i:�
frhl���9NŸ�.��%��)�X��f�ZܟAp��~ģ�DEkY��-��aA��$�ɂ>�K��
��-�p��j�|�	t6�p�]���8=��t�A ��r ��/��V�N��|^�-��9�;�,� �#T���:��B���㓧K@��*�:����#���3u�`�x҆��I��ҽ�L�Z���(����F�ںe����Z��d����j�1�u�.O"֝�bqlw���nGf>Ƨ�:�U��Wn�}��J�b��EV���i��cQ���K�1�QQU�M2�(�HU ��\����V_�ƟV��5Ȃ-\rFX��=�c�B��d���r��j�b��3TtF�?uD
�@�&1\J����f�M�6i��q|Y��)��$��������f��r��$�����? �֝�	�8w�R�������D� H������)�-��_�/��ڹq)Y�13l4�r�8�����EMd�Z�f���U���#��v��JPM����ہ3狉ӺDJc�p1M2q<茡����T��Z�-�3B�����.�6�#\(P��l۠����݌C�G�3*�C����Q,��&#�e���[k���O�2�vqt�:s�C�\��B�@�Ex-b�*Jk�?Z�R�'���$/L Ÿ=$jK���)b0P�Tk�w������8��JH#$�}�΅u�r:4HA�Z�����/�1�Tf����a��.���s?���%��罜��Uq{.>t�W3���#Bj�u���ҧ��M#d��p�e�c��!�Y�VmS���BS��J�g�Lqu8p9����q�*�˨~Z��E�o&a*�q�徼+����8G�R��^���c�����(0���-d3vF������B�k~��_7e`מc����aœ��q�x�\_�!x�N�/�,�����*n�]4!k���2�)��೵���g�@XW+�:.f�1����*��Z�Oy�H'&�u��U$��'|��".HG��K�s���1��o�;�
�_����k�s'��MȱW��Qb=~�	Q��}��x���6��ݧ��bI�S�F�q��At�I�F��b����� ��#�����GE�MA�_G s��3lbE��?iq�]�C�n�uI�5�t]N��)��I �7���!R6T&�s�a�7ZDPՈ*ڎ���*��U��чY�ږJ�y��{���\h�T�"o�Q����߱�`�7�m8H�X��}[P�H՗��L�������q��B�e���Ec��jJ*!��1�h����㸗-V�'KU��(CC���ٔ�W�J����"�I�,fӁ?�f�,Uf�#N�4�l5��%t�z�bŔ*�!W"WXG��e7U%�{����j�0n_��T��?��^&��>DT$Y�����, ���j1G*»p�5���J�S;F�F0��j�����1{�M�G:;w<HD�f#�IMr��х�תJr�'&���z�k�/?�r68��軡72g6����[�:y�x�5�Q�[3�NI����`�7}�yeH#�W�mN~���w�����C�@�4��v�:�
m��4� 7�n��)d��#�{�J�Fϱ���$K����8��r��4��m�����}A�T��JP�f�Jf3#�c�;y�`y$���#�P����Z�����3Hͧ�H� 	�t�gcm�'|hu�虊�on�2���{\&�Z�M�rO�727�8IxgQ\��-ܮw���c	�T@��e�I�oŵ4Dԛ����S�i�ys ��03�N��;ǀE��������<����	��@^�|�.9`�D�)�4�N
���OT_�̢�3w�x�������v<Ւ X���}�VJ \}΅������U�!�x�d�L����]ϴ%
�2c%�d��+�z/�$p���A�wx�,f�߹Q��Fs}����D[���V�MH
o��|&���n ���g�ç�)e�x����=H	�q5p��dlr��W#%�W�tŸΤ��G5���.\r�����"|6QIK���Rb�����g�1��$����I��T|аwR����l�s�y��g�'�6J��aN���y�?˨ x_!&�e0���T8�����ʩ+�P�H�C��q�e�S!�g6�|����V3>{�5+֮�O�k+W��
������d��O�sp�T���/I9z�f�@ۏ����>��t��˜����x{�����ey�z��c3�ϔ5�{�ӎb7�V��CK���5u����U���dGo�Z�l�.�(�\r�`�aV�a�y��&(��&�?�Ǒ�p�����T�ѓ���"�"��#��!��,����	G�eGx��^\:����W�$Ax,��wX^��t^V5�u�ܺ:��k�~C���ɘ*��d��X�!&2���t�.�������Ϯ(U�.I3���/���T�(�y�C# �k������q����NC��0�|�I�����/n�c�D ��7��э;��-cjr?u*�A�>M��Z#P��_��=���0�n/�	x���&�Ԑd�R=W@�^��WYn����F%�!!��E�Z��	���s���@o"6�;q�u1��S�޴��_�>��И��I#-�K~~
(���Ѷ�|-*a�ά���vT�?{�<PLSM�YTAe$q�JTZ��UU�TU�q�*��3��� �FI�z���T��N�Y��+�*[K'3oɬ�Dav'l5ٟ����1mc���_�Ȁ~x����,ة>�����R6V��Ճ��v���-���c��86�+��$����.�5��S����H�EL6{�r���4�b�	��I��2�#���&*D�VZ�Rv<�}[��3hR�D�#ې@�.��^D��6<Ǥ>iU���;ǰ������dt|m��9T>j� ��rR�t̬ ���+Q0z^K[,C�^�#���`��~�*��,�'�G/ۤL4��	 {!̴�b7�mZ�������}�&)׊��A�����DH�1�m�/���S��S[v�rTۛ�w�C�2�u:���1*��i���jpE�Qc�b�r�.��X��^��,�9�O,�L$��pF��Ϳ�b	���^In��Z�j�>�չ]�Z�c�q�v d��! ��v�����(��7 iZ������24䫂�H*r�bhj�K��#)Z��B�g��%����9���+�p����Le��U�`�s[���>��YX��ia��_��,��p��L�cLO$�͟�)�
hz^�2��քcHYV�(���,;�����0�Y��9��YAֱ�`����xzK7�?Z��U�z�JU�qE0�CV���������%|S:�7%�O/���Q��?���8�nwUnd�ֱ��k�T,��}�#�6�h݃��vk�!1|���Q�Cn��L����z�)bZG�.�\t(<<q{�x��bF�c�= @k����0	4/�8�ǣ�
�P� �ijM�#�7榹��N�6@��3��=Ȥ@]EY\����H0�]���L�,��e�O�9�?����筶�EH�(����iofK�����?w�/(��KQ<��V ��9e��ݦ��:�
�D��Km����٤��Ey����r-�5@���㼓�����D-G_;�J6���b �C���#MP��vW>���Q��KZp$bm���1�]�e�R?����(��yWM,Hwtj��3�Ɏ]�Ĝ�n9X��N9Y���u���6I�?��P���1Bz��b��5��/*ǟ�>4����߸�m�i7/�E�~�P�M�Р�6���%���ry6VXk�\�)�t��sP-m�����[��YX� �息���;��d`�L1�N��i�Z
Y�BY��ω���P�ݸ�6ͮ�����a���% [�V8Y��/r-�����h%O����\�Va3���dB�4����-ώ�|fL諃��e�����y���]��oW��bB��j��pu����h�~ˋ�O��.��,GI�cK�픧��������;(�FH q��E����\����d�*�Vd�s�O7��/�`�d�}9�d�~�h������ _%l�o�p��BK�� �:��'�`��K�@�:oM������D0�My�}j:P|&E���V��;y C9 (�cShƖ�3��9� ���a������<��0�Og�W���D��_�n'I��i!��4û��?!S��R��=J�c�u;�*��,�iw�[�ߓ:���E:a�\z�{��3���(�iA��F�!�Wwc-��=�2�{���k�uՀoݟ4ZF�,����-p�����k�~���[��X��y����sj<�ؾi�\�zؾG湢H�hJ|�&B�]�� UR�ްn��e�;ɔ{3��1b��$��81�@���d)TW�5��dc>��D�P�\f��u�����t˴Ui �Y�`r�l� �SRG˖=��׹�Q�$�uSݣ��&����~�7͓x�zLH_���� �=W:�4?�l����A���_B�UPg*�nh?ڎ���	�Ʈ���bt���"�U�a�/gs�4��aο��_��F�Dm��
Y�}H��oIo��@I�ZpFL~���䐔�����(�f�k�{Ɔ�!W�.��`���el�L2d=PL��ʮ1���}�R�zӎcH�Z�c�����T�j[DI�g7u�& /�@"	���B��ax�e��TG2��m��� L��h;�����)�i�d�s�Ů��M�ǻG)ش��+��6�A�����Wr�d�0*0Ԍ-VH��̴��2� ��ԵN���í>(�*��q��"Xm�D� ���Y'����9�w��?�8o]%E�GH |R��YE�=kx���>� ��e)�>2�����xg�n�g��'��� =gߺu��;U�2Y]�VW_�gW��Su�;�	c�J��%U�|�%��E�[�u!�U��Ł���v�:Jޟ�J:'ć�f�=u�5�{m*�c�V|�*(�כ��X>\$����8*��h��������A��߅��)>�9�{t��N3�(�s_c.�ɣ� Ԯ�SHC`� ��=��*	
ɦ�Ს���}�E)��Β����R�RuHb	��������Kx�C	�s�)�vY��ٮ"��D�EQ��_)�j���e�L !�Ӹ`*��__�@aQ�ɘ.R����@&�,y׽/�fF��w<[v��ƒ�)?KÄ���)��Xgv([�\	�L�"�9�s�%bk�u���ڗKÂ�KH�Ci���?b~�^'לD|!���f_�dt�=5�H����R��p1A�����mQM���ˆ�.V�@�9�a�A����>��b%��<��I(�U�8_&�7g��U�dZ�µy�g�%)���P0i��U�io�I�nf�!w�3��+O�H�v<����:��C�W�NZ��` ��`筃R�,";i�*Ud Ĝp�=�bϚ��}HԿ!F��E
�%�*�=��@}�״�tM.�������T�g���&�;Y�i7��CgqT,*0�q���:�͇��������&��;�5��;_�թ	#�c���%& MN!{^�-�}-��V(��E�v:|��t��R\�Cy�W�kN_����]9d�CDoH@����]h���3�ʻ=�SVw�ކ��u������s����y��x�V7Q�.��+?��NH�W}?�㨬��O���~�m��)$�"]O�,�=X2��_ԓt�ᶟ�3nY��N���{�݉Kأ���
\R�j���������<�;��*ޥ�Nt�>=Q�V����:U���y^0h[�TG��B"E��<��rH׾�d_�x���`�3Fd�;�{_���ݨV�������O���_�'�V4DP�E��-C��܈����q�6b��ov5������E>Ft�~�|+���n�]{�m�������{ი�C�c(s�WX�|>.1r|�W�f���Q�j��T��(;��̍c����NZ������_��j�~t�"3�iv��uS]h4�5���2n�|h�`;z�Y�Ζ�Y���d��8�K�g*�h+�s07W�+!73�ˤ�$�N!	V�f�r�$�����Y��
���e�X��h��iM)B��䧪��
@^Ks,���,}&�~^%�|T�!f�Ո|=#�w��]�X �.o+.�h_�񨩮.[;�yT|�.<�؍%���w�rR���)u�ب}:�\��h�a$�ݵ��4`�х��Xe'	�9���� "ZFz�@O��9�S�4����vpvL�m�8��t�TQ�1� y���(�b]9�鰊]�xA,��@��`V""�o�Gx�Ye*<rnӘ?�S����g�&�H��/�%`N{hߜ�!,����(#���rig(�KV�R�O�ڇƆL%G2�J=�/�t�Ǵt�aJy����1�)I���~1����t38�2L���GbL1�I���O��ƥ�#aF*�SSd�k+8���{�/�=�/��E@=
X��W�צ���Ҭ�����;3���Ȱ^9�D��}=\�ZI���V}�4����s���O��҂gR@w_J�>��p���eM(�x ٪8�it�曷Z��lr�4k�n>I2���J/��/o\��β�'�����^��/��\��2�N�16_����_b�F��z��f,�5!�=3�$7s�i/+���쯋~[o��0$�U�&e�uL��1&E��D��uRJœ%��4� ���A�	�f�A(6SK���'�N=����:��o

��ԣ��0B�m�B�^R�3���|b�I�����l�c�k�$����^|B�A�el��d$��Ւr�`�V>���qVmD�&"������)��>��h�x��p_�)b�٣ڕX�W~���ȕx������@@�-�%���>�T�����[z��k¢�P�5!����u�^4[-�0J��;�w�h8���?�%R�"ǋ���-��r��
#�X-�OJ��p���r��J�]	r���.���6��[h�anUd ���ħ���>x�)�4�LF�%.f�Y����^h��r�����7����k�)����MnM��C< ��q�ӕ�)���U䂏�aM�_o��j�V��'�'�~�+���Ჸ��N�N����g���v�k~�\^�m�x�����O���9:��m�;�P5k���Km6�?f�e���2�?4ns��@�� �p��{��⎜D�HE��՛�x>2�1��a��^^�i���އ�8��E���"�Ѧ�U'N��C
l8Gs[Gb�V�^�	%q�Q#SEq��;�7Z>�K��9ǚ0�L���-� _g�	��P,�2~��I�� +��/+8��q�ʀw ��1`v�?�L�3U�ŝ]Sn�㶪q�_��Iw�����DD�M?N�:��	�ޡ/I �8E�B� L$Gt<�(8��,��1�/��b�[��u~�]㺙��gs��_s��I�V-��
�b�"JnI�!�*i&�����"��oB6#��5ʀ8��2�%���֞�eթ��z}).�7ڠ���生Ô�G�8��Ȟ:_@��7��%Y1S2��'�'�)
7ہ�C����*?�%g����z�*q]N
��2~Lrd��1C�@8l3�u�����R��i��G*�'�vnF��$�o3���� �qM&�FK3]�I
�����UvX+!g� =��ϲ��6�M"3w(��3���dW98P)`c{If�-6R���]M��ag��ՠk�bH�	��LR�Eۮ\����"8�|D��A�����a�>����zzp\OqBd���x�qY6ԗI�r.��e��l�c��+=Z>�W��[Keҫ�w�?�R��<�l�Q��S@��/��� _���q��ȟQ�81�Q�9Ń̗�9\+-%���Z��a�:�����I��b^�	A�G��,�}<Q<�{���'-����oy�⨦?�>:qu��ۮ�3�ns@j�nK�
�X
iz�G�Itl|�iM�;_@Y|!�D 0
+�EL�&�+q�Q��)�m�%J]���!�:7�u�M���8h0h��ace~�Ʌ1�;��=_�*�P�➥a]�AE��b��+݃�k�`�/̧�[C���lA ��@�:��SfA��c��y�vV=QBr����<.e���Nb��B����[�2f���5\A)�X�yɴ$���s����ԋ^m����2NZXԋ^7����=~.�����?A��;4zy:�7E��H^1f_�©,�*��x�z�7-B�G[��̺���5�9�����1F�����X.��T�piU���4����9JqF%�zh��'=�`�>���y�~B�i!<]���@j�?���K�F}n�:B�WU`����<�C�Y�._�f�a���{Ǳ�e�B02�G��rG���C�7��V��m��z�>8��Yjg�bX`F��t��.
��rH6��^�X��?�R��\�D˭~3��h�q�"����^�
]Ȃ�Cnr� ��K ��8���qKI��!��P�<'.����*ˮ����
��-K�sYM�5����|�6�.��9�RK9�$zs�!,��D6��0�'�J�}��Hq	��+.�Vz}�i%�6T"�=�Ҭ��EXi�&K3t�h����y���Q k�n����E�e�YYL�ɐg��%�d-۾��!TZl�b�3��+���9#��WC�E�yv;�=zɣ�3�K9��|�T����J���G�Ђ��t�E���̂Cљ�gB���fS�!���5�6ޔ��ĥ�>�nF�V�
��q���\>��^�-\x3��7��Sҭ�8��M�*�h������~�WE*�t-RU�0�I��}��IR�g|ϹI7G��o��U��[�����!k�h
D!,��'QMVF�!�H��g�SZ�g+4����t�M�������V�q?4��Z���Lӛ�Ӄ��	�9B�=������aad�� ��� i�����w)�3�9�����x�'2�j��N��2v��+ Jw����ur�y���s��Է�x��w�C�$<$}�)���/�02H���J�~�2��\u^����Ơ��̂s[ݭ~�#|6�5����7*i*��Y��,�Y��V���7�?3~
�B^�/��d�(���%4����Wb�PgyhV'�h���e�F��%AL�q�����)r��v�:��ëעذ�,��~+�zw��@�\�XR�k�]�j�����B���T�1����i���6�gy�֌s��s�
��SgSfux�`P�Q�3O��]	>�U��979[>�?��K\����ГA[�`*p6n��8o�q�x��^Al��/��u��PG���W�?=����#?aꢖ�>MUo!bƎ�&2|��pY�ȥ���UE�_xUT�PX&Y�c��ۮ���S� ��ϲ'~�����Rp��-<Ÿ�}4��N�Ns(G�ݛk��ZJS�u:*�Cnh6�	J.��E�9G������b���i�$�!
�U�^2~��d���]���#�O,�?+2�*nN��L#�/���z���\h�'��G��W�g8��MpR�F�������4>���O	�1�x��K�#��úlkg�+�m�[���U��� "4�J��Tr���Y8a�k� ٭}7�<�F.���>m�b�5#�uu�Q�f�$��+�����6v6����*%����|��8R������y�\)2�&�@�"$��zk���a�f�+�X%�ܦ3QwaG������{qY����!�%��ק�:��%<�".�'�+�e�[,$�W�".�v5���2F�;逈 �n�1�4P�r�~���ɵd�������}ʥ�I��*���y6��DC�I��*H��~:��)�m�'"��!8�.?�瘸�Z�X|�<X=ZR��I�d���zO���C)ȏ-s��,FvTis�Q¦�����[D��#��oE��q��e�� �1�Ս�K�H�0���.x؏�#5ڱ����ly̒��}Pn�<��B&0U�� j�� �l-��>j�ϙ���0~Ȼ����6b����}瑑�[(��1_G��xM��R(	�Y5�}Y5�\DV��Z�HA�����w�H�a��{��4و�b�#��}�ef&�e �Ї�8�L ��Cr�I<�+�p�M�h�WY���ҙ1�OB+4	?w}�9��7��_j����Z�>�u4�+��� _����Y�z���w���6�5�f���ڬH�ia�����j���z�R�ۭM���ɛH|Y��?=[� �Y����O��}��l#��	��P��d�����~��gu�Ks��.�"�/=})ݿ�^����˷����R��/�_}�.++��V�66���*�`�
u��p��Ķ��v�`R���.���!�R�jgbd]g��z�}�\��5�5�"JH8������%���(������	���,kM`ʼY���.1�.p�i)��b�	Ј������'�1
n���Xץ?onn}s���3��s.`�<r��}����&�s�7�"��nL�}+�|�b-M��֊Ya|&f7�=���n��l�7!.N�����/Z#ޟ���g�כz�v�K^-]��5'e^��JJ�o g��0̀ ����<%�m��=v�<�mç�S$d㎭��0?3��Ǟ���aU���EpB'�sC��CX;�f�{}�u7����;D�q�P\�Z����D`Q2u]i��
jA�KY�,���"�g�}lv<E��F�418"�;��@5��k���i[��˭��%�S{~���s���ʛg��܈:T�����3� ���&���i)�Ț��Ad<@F�g�2Ջl����+�84���1��X��ה<Ș�{�)f�r����8Ùu&��Q�2q�Gz�l�&��rm����t3a�/V�z2s=w�������u,c��%��~�VR�����(|No����~U�\� �(
���$����_�+��0.�[¤=�C���ca����)�G���ڳZr��s�O���@lb�f[u�������!_[�3l|���b׿�ݨ[U��7\�vuIN�*�Tկ��yC0�k�MMr29�H	YT��f��߂D���S4ªJ]@�9�G0%S=bG���k�8�O��� �@HD��\��kK2��#q B֥��^o�� �r�F)T��5c�����~s��������8�W:��&��ZG�x�;҇��J�0�C�7�]����g@Cid�Z�GxƧ��W����p�8����m�$�s�Ӭ�?�e]ѐO!q��#C*|���~3$D�`}Ibw*����2^}
��Dm�h�5����2т��*8��L�v$�����;f�31�B��V[}�z~��Y,1�"��-��d3�p�Yr'~���r�`LT����A�r�?�G@:ÑAiX	#\ �JD�ӧ��=��B��\up�ug�����q�������o�{���P��L4"������x;bQ�p1���˔H��ҫs۪�=A
/ߟȮ2t7$�6�Q׷b��gkaXfv��_5��
�cdN�+�H������+�b����Փ]l��D�g@+�*P�/s|ŧX�f!��9�	�Z����~��Ǽ���L�>�A���DIQ������w`���U�ݘd�UJo��U���A`��<�X���Y�1N��RT�)�z�܀�m
�NƄ�>��:���Q��)�abz�'�&Y���(��&H���W0�j����bX����x����г��c`_Dθ/Ǵ x\k�אU�J��[P$�/	��?Pr�l�A֍|� ���I�'��R8e�O���I��%Z��Z>[���>@G5w�}�u]v�-g��K~S�)q^�q/Tnu6��lCh%B�30<�����@؉�S�7U"6�*�"�M�����sZ�|T!�"Q'ݎ�>N��|7�9Y��O��u�{{�w���v��"H��\9H�k;�W�䀌�Gы��?����{�������ac�ޏ��H��
&�0O!$#��C���4� �4'v��MB�6�Y䯠@�u���J$��/0/�}�����"N�1T�
���F�M�s&��D�a]K�����g!����Z��{,-��ޒ�|_�95o�k��c[�fضR��zQ�*����/*#	��~�-�s�_a#$l�<��!����%�t��|T� d�}5�F��J(�䙱Ѓ��}g�St���
'Y���}��a�l���m�m�@����d���$�wp/�y�6*��X�_p�V��1�Y��d�\砭��,�9�׃���J�x�\
���F3��|W������ú!icI��F|��Y�H[A���!�o��R~o~Y�Ej�W.J'+� .W��ɒM/�#�]��FH���dO ��l�Ʋ�<?܂G�kѧ��e~���i"4r�A��%�4{��h�I�����ZY�<"b����M�����Qg� �|���7�����+SÓⴢ��WJ�1J��}��zd�[��������䩛�> t�-�(w �`�[�'�|���V����1+�S�b7]^��}�x�s;���}݈4d�1p!Vh,v����E��`i��{�&��(N���{E�w�O|�Di�L��)sԉ)"A� ��	�Ϸk�������O�S�h��}��G^en�]��3�#"���`0An�E��/��\�#F_(�ᱢ��0�"u a/Q)�}
[�c��fy	v��%o���Z�kRJ!N�`,��Ӡ��2�l�V�� �Ed@F)$��%��E-��8(�@��w�i����
���(��5�k �En�@�7Oi]����9z���1k��"������8d�_}A;���O���D��:A�7lߡ��	|��6(���D�T5Qހ"�莛!���%7�a~n�Te�$�@�Wdh&T=],�$��Z�;��~ͬ��#><��!-кb�E=�V�3��C�������0z�#~3 �JLW_ͷ6�l6�,[���w�L�k:��G��u~�*Wo�"�h+8��iѐ ��q���z��r;PV�OH�gr����D"�v
�Ù��\�R��;���H8"�;������tm/��F�l�����6�4i&�ϑb�I{ *����v��|�'��9��~9�A�rꤸ(�T�K��
K�q*="XS[4�߶ چ�\�/���T|ɿ�m����7O��O��~��0G�����\˛ӯ(��=�{�b��Ǧ��cn��|��k��V�B�����M��݆�H,������*pi�D����#�?�C�:�?��|��ѡC�h��tM:'��ۍ�#��l��~�{�o����wro�����G.j/��/qPȍ��4X��W6��dV@I��礂��w�ɡ��~���;�vҨh���`h���>E[X�ֺfr{���\��ji)*l}�����2���~�@Y��-~�}oN����k���q��<Js�f�;�V�"8�z���^+��ϫ޸d �۳�4�@�	qS��;40������u��c[3��[����xG�����疪`	E���C��c��bF�O��t&ֶ14O�~S?�ym~m���6�so4���΅	Vҋk�. JA*wذ��J�5�'
k���;�fMzx=�/vƽ�}D��nBwH�֝x5-��N�ZVgܤ��"r&'� �U�T�Nf�V���T�q�Ǣ�$h�S@*8��n�l��kDM�@��dU��ao6���0�B�������/Aoķ����j�i�d�1�*�:sK�a� uju*%(�5�����]���f��3��	���WX���/�&@-����CT���1�օ��aW �e�M#;F�$P�z�T����4ES�60k��U���j_^�ʝŖ/��ڈX�墫^� @��)�rJ�om�՞ �j�/��iM�{b�lȏ5]��@�������2~O0��F�Iv5�W�+�rE�X8-?/��Jyy�O�=�]�~U`<
WN��87��<M]���+3+���kLiC�I�;-���,��J�q�Y ̐�$�ck'��ZHw1�J��/�����9h�S`��m���ra\_���(�����4�q�J��
�1�����=`EC�!��Bo��������d��}�����C��?k&bG2e�r��4��	��e��0�kQ���J����L��� kޭ�=�\���k��#��e\[�DF����.<�3a���N��ie��F������n�1,��%�L|l}�%?�竧�<5�R�ZQA�iH��˝��O��*P���Dͺ�9��+�l�HM<�Oz�-���
aF%�8���.�޴A~|@Y���S���z>&�E���8�H��_\iE��: e�N���S���
���m�ߏ�����Cb�4}��E弸�Ad��O�3�Gq]'S0�P��G����Ia�nξ�<�����%Л����mHH���F^8MXљd�'fz�oR�z�u�r��˓�:���t���?C�I��D�R��lZV)��3����r���Fs$0��������<��)t��~~0���L~6���(�gl����q�FJ�lW��/���#gX��Ϝ�C��dzc�7��8���������ۄ0d�V��=�"�ѧ��.wR5t�}���I��:s��&z�#u�F�F{�5x�@���kV��|�]S7Ҋ��ʟ-MD������ӥ{�����\�6��������rz�r}��o�K��8"��^���K����'哝|H���uL@~;
�/��Z��p��<	Ē��K2�thV�.7�d=5�碋̅�Gp8k���1K"j�T?�#�{v�������@�萏l,!�!����D���B/	�^�<���sP�W��㸫
F�<���"+���:O�Y��2�蟭'o�M�mvwڀjc��
Y,RS�%��8a[�Ε'��9H�����)�����5�k�ò{"�	��C�C��2���ӏ�-n;��cl�)��h�{��ǭ-���q�?�0N����m! �9G�9F��o�cO��4��z�Nm�z��qZ�ۢ/У�������l�m%O7�XH�fM#�/�{�e��4�ªE���-S�}�il��>�-��k���ě��V ���C�Bz5^M��ه��'�(����Υo��0ې�1-jD���9'%6�fg����;���eݿ%T#ᡁ�ľ��2�����@�>Q��-%�� �O��.Kz�d#�0c��&������,��a�i�I,y�	w���,�y[Cb��l�+�וBu4��]Z[�Ԇ<(𴏯N���Mh���&q���T���5��W�����x9ȕP�m��v�-�����������a�>*.W-"��ɬ:ݭ�$�HIS�˞�b?�`�<K����9��'��m�5|������%)4�u�Y����^K�ްC��Үc6D��{���sP�
�qy)0z-,~=�>P���*�*7���3_��.p}wSd�X�>�U'���>8,����c.�'2��B�1��2�wo����^���k��G��n��C��D~l� He�-�V�8�:r@U7�k�єuf�b��	��C��)������/:����&��^�G�8�U��J.����~����ǟ�3��XJ~���Ǡ�� �`��GΦ�vuW����Q���H�n0��Obq4��A����[x�OTpoIt�S�}s�g&!]:eE�:{4�j[�!���\�mԢ�Q��K$lIg�2���=~W�~k'6q�Y!@fu4�)�m���ȩ[��7t�0&{�[�x4N�y�C"�gF��Q_��B�=52���#F��WQ�5����Ƚୀq���p�+>e�-�N���Z�P�ΰ;g�����.�3�&�<>�2���Ah|��cy�:�N�q�~��d���B8��(ߞ�>��O�i�q����즂(o���s��f�3�a�m �#ks��ܜ��*漣�WzfL��F��VK��nw��4M��q��{����������tX/��Lp�˒aK$����~���Z�Dn�5X1�|N;g�m3Z���)�#����s`����:ߚ{s��$˿Ә�dO}P*�hf���c"��{d��*�<�%x{�����S<�U���^&�3�Я��M��2�1��ÿ��ƵM���7eo�T�d��M��Y��y�vҤ����G_���v��p�x$�z��tB��G�z�p��ԧ�R�y�*�JO����|2ѷ<��\�=h����r����Gk�e�N�O��n��Pi�1��������շ�vkr�e$��F�D����^��P�����Qb�^B��ˡr�F}�ݬ���K8�=�*7��ǹ�
�u��R�]e7���Ѭ�'͠�+�so�"�Ǖ�Y�R;Dt���ߦp�<�At�+v�
��Ɩ�ǁ��뇢�����<!.m��!'u���(7� /UT��Fr�=!�M���,�sl_8B�y���ur'�ـ��~׉q;�0ޢ���y��rչgH�����?)Eb��!��Vh��|��P�Q W��,������T\�l�u	1���;IR0oGV�}��E)_���0/\�l0�\�;����v�O]o����w��4�Qt��'D�����'�tD��{6=����[��bh
(2��|��0	�Ai����+B�%{ݨ�m�r�g���[�f�ˮ�Ny�6р�_�͐䬘�{p�әX����B���sP%QQ�qH` ���C�p[��j̖�����y(�޸i��@���Py�[4���	1.��D�ᘍ��?�0֑n�γ��-n#�4~܆��,2�أs88X�4NT�B��L	��R6#d��8�hG��8����xz�l��~�9"�����:3Pu�N�\P�ȭ�d�p�|渋w�o��p�g��{m/��L K��O�vE����b¦�暊O�8�>SX�_`�s �}���G3!Đ:��"��?Q�&��8���֒?&��Ƞ&pT)7�֖(*o`?��a�hq�=�G1�	z`[T��Ƭ ��8��d��`)�,҃��1)��^�qto�����\���� ��#�^�cIz������³�w����A�J�����9]YN��G&߸��6��rD.%?�0���������t�V����}�E���>/�����)0�Y��᭰*��!��~�q�k9���i�(	&0�x1�QL
}��xV���S�ԯ��"�|�ם(��Hp_�S?4U����9�1X�6������-�ge�{7�\O
���*|� oy\���S�����Ֆ-�k�)~��6�i��~TK^,�d�m��5��]uN��FJR6a�&�ʘM?��! ��m~�����\)K��(�N�Qv5�&�,����m���zVL!?𕫚S;��a��5����z0��ґ�����Xy��y��]���l������q��#���@!���l�?��`��:v��v��QED����3�z��aH�ds� ��[2�'��$�����F{7��΄���ý����7���Z��*�L��M&���U���[�ߖN�"�Z���z�:�Od�7�>�&ӓ�z�ESY�g.M
#>� &S8�:�ȕ�Zҕ���a���m�تV��lR:�/8�x��5
�U�ݔQ����htû����m)��r��:��WW9��;�����G0h�3�D��}�z�A��=�cv	OMor�*����u*�5d́��b,ޣt!eU�jWX[�ŲC���#�������T��1"��k�E��)i�Z;,|ͤ�WԖiK�7 � K��5F��0���0fA;sA,�\��e��`;���
���N4I�9`ྴˉO���}�v�v~�Ʊi��Bj��'��|�ӓ�w��#Vt��YX�3�p#
|J՝C(^����Gɉe��<�o�\Z05��:f�Jft;��yz�u�r�8аĊ7�b<��"���<}97��2Ӟ�}9���%�����"t���X1+E�D��M|��R�9�((�rbZ\+�$�էz��afH�@z0:11�9jJ�^������F!v��jlS�<�����H��(�[2 sk߾f�X���i�
S�)�-�橣bpO�8m��:�����B����|�B�š������c�`��T)�5vȂ��M��� p�Y�M�6�O�&����b����F4�x*A}{�ϡ��)�D�Q���"�BhH��d�����K��/����W�(�0���D�I��o�����2Ʌ9����B(��*,z�x���lںEC�q Cp1��4�C�O鵪P�JY�ac�G���}ߕ�c��2I�\w	/���/�zGDg���1�yA��a`?0=�V��Cm]���Z}1TlH2K1GWM�䯏��0�֝�F��l��+Fn/:jL�~Mh^��#��7���\��X�
������I��x%�8�$&k�0����V�^d_�<מ[�:R�]zC�|�D���Tpuo�h2��׻X�O�ɵ�qGRU�l_
�~|�1_Mu�Ls��M}V���Rc��L�{aq�ʪǧG(�}����h�OL�pȱ}T���a�ݿi9d�v9p�|n<��2I��6PU��H����N՘'���|.��\k"���@9RJ���-�{��Sl�7Om�i�d�s�R��ٝ*�[Ѩ�c�]u�͟T����M	���c���H�I�o�0� �_q�?��=�'�{x�g���I�!�����}kLh��I�n�/q�4,4� `���q3 �I��d��Wp��� �*Ò�}gD��Y� ���}�LJ�>��]~��Sٝ,cG��5���������K�ǒ�NE����n'�7R�=�H��`̰t� 1�X��I����/�@����������8Oe �ܚ��VK��7����uX�e36���azϟ8iPw_Ty��í�Ɖ(�����7ٻ�Wm❹���@��q������}ܼ�����V�yd7V+}��9��&F�Ya-���A�La�&�Q�Z�;�}�~�����z�*�&r�qi��"��-��jrhd��Z�d���/I����W���nDx�����c��dJiD��	�g�����͓l�a��T�Y�gz+:b����Y�A�f����x�3�S�2{ 6M�z���}�f�鬶�T�L�K�Qw$�qQPԁצ�`�ex�ڤ�@��$��� ���
�I�GHd��uw�2�d)ы����_,
���Q+C#!Lg^c�T��6;y.h�ohE�<n����>��)�X3CD�-9:$s
��:%��ȭR%���Eb^B$g��C�VD<� UMM!~��u!>��ʚ���lc��%����w�'��CJ$��]�2��(���_�mS͠�r�\ۊc>,�!�ܫU3e�܃`k)>1���X2��V>-D�$n�������ѐ��s.�>��UZƤ�4��.��,;��Zt�w���d�N �逊(�k���ދt��*�,I�� z�H:�p���o��t��]�w����.�Մ�n�TC�^�֩���vt���!A���w��`
��%�� '��X+��A0��C*C��r��o}��(�ǻ�n�U>6���U ��A��8a��&��9��Z[>sU{p�l���q	���[X��"���Q�Z(n��jѸ���6��=���F����e;A���<��n��OОr�DF{[��;2��e�ꨂ��K�cY��i��C֭Z�![俥�Oq�ω<7IJ_n>&��교b"�|b�ҧG�����n]�)���i�������I蕮����&���{��	��z�Ȕr��iީcU��'o;������χ��q�E�9}Djw�4w�^�H� >z�Y�����s!Z~���<�}Sa��Æ ��=�3
��hOIc��2�i�p��@
o[yU8�FT�q��p��E3��-ʄ����/r�)�T�����[��ʑ��z�`��9n}|4�2o��7��M[�b�8)�~�z	ň�#���ja�<�/N�G�j���RZ<vZ����A�s	�]�
N��Dm���Hn�*89R�0�+�x���r*7��d5i�%��?�i�<v��E!�T��˩wv�캭�<E�]�b�]�#�k���{	l��a�Ƅͩ�`չ|�CX���	��Ά����nOB��
�$B��L�S���p��n|=ob����K��st5��>c������v�	���T@�Y�@�4bw>ޑ�]��	�>TB0��}���lF]�-2g��E8�	cWO��T�?�QqL��
,c
9zS%;2��e�&�n,��b��m�*3DMvac3cQs�����*�'P�E�|���$����jK����q������S�D�:�������'"�	th遮;]X:���cXrV��c{y��ϐi�����/d�.'��7�}_7�D�2���l������N϶���J�w4ƒ�
�a�v���B��{"��wup��{W���M1�2Z���k�z-��b�a�|�MB$8C�[�jL�N;�
�M��K�QӤص\U�*���c��ȟHN������^܃�[���p��~�2\�e3׬h�zu�k�u9����8�(��^n�J��3,�0e��[��x�~�T�����3�\�Gנ{ j���ʐ�-�ƿG�V�|�>n�v�u��X@�JeΖ�*�s^!|L�O9G1�&�q�OD���8����k�P���|?Z٠*�J]�6��Zc�Y�.���r��<��
���(�/�H����˘�3�i��Eu|CZp�.l ��$�����v<|�������m�s�&�Wނ��;`��4����.����OǘT �@��Y>��4`�va�����8�Tc��^�p�UD�j��r��.u5��a��&[k?=�9Ε/oO~L��M�#��j~&_�/����U�Ů�����<�ى��օ�cr��Z�aBm�[
Ǘv�<
�=/�����H�)|�9դ�%���'^�#Sm��2l-G�r�L,�K�aO�����9�^�f�����i�����2ڏd��ݶ�:r���,�j��ƲP}��o�y]jj�0-�*���P����$�_eu0��q�+�����L6��*}�f����Y��l��B��lXc��J|�g���2�mq��%R��퐭���z�q��6b����ҍ�"@@���u��c�B��ȗ6D��ɛB����◾��W���O&��Tq���7w��#wvW��w�豮R����js@�
�q��< �&�YT�j+:�v��5�Z��݁��7�^��x*��K|>(�B�������m=�8k�B�-����ڒջ���������W����K!����u����+��v�?�8�jOpZt��k��N����$��������Re���Kѝ��=�������>U�wة`:s�u+�k���]���q�� K�k�;�jнޱ�x=uG�)�/�'t��^�f��џۚ��ͷn)��ۿv�����}/-�r���f��C񲗣x�u5
�
2_��M{j����zy	 sS,4�� ��h�ڠl�����P�"!$����宺Er�!C��찳�.,��}�IY/��0X��/�O�k��ץ�c(uM�QIJ��$z��z��B��d̸�b`*���;Ֆh��fk!�V� �8�D���j^.�{T+��c�J�1`��v�������� ���s9o�e���v�����I��T�K5ݔG�r�
�Q��|7����F���-حй&����UmSR���o}��E�˘]�ȧ
`XI/��d�#�'v���Ug�P�Q�{h�7�m]c|I�w�$s�z�Q��P =��Vw�@럅^EfQ2���p���f�v�PW�Rܷ���~ې�lz������TX��7�[͸��`���`U��	���)B�E��*Rm:Fe���O��>j/k���hHʆx�{�6��EG��'ď|8��Db?�>��^����d��Z9����; N��&a�����	H��Ʉ*��L��VF֗N<�82�}�U\+�Ԇ�{��!c�dz8�LE�Y����^l S��[
�>nlT��نG�8:�t���bR�Pۣ�&�y�F�@^������	&��t<�_L0#B��(G�эB�?R/T�Eb}��2�����Ӣtm��z�aͿ ���oj��W1T���Ȏ�W�"h��1���L�H!SȖ�I�^ROvg�f#�cil/��J����9�y���l�e�h��wJ���Z��[9�U�&�s��[��&�κ�ok?-������0#J�/R[�s�����EY|ڶ��pz���]�/�!�F��݃�/V�v���R�|��������BWA=��߻{�a�T���!ͷ4�Rls��*���`%�4�j�4�5�����|������	�3�ߌ�?WX�I�9u�?��K%�T��i�cx���ݛ� =z��.�8�I��6[�'3�K��C^2�	R�#�J)�����.I��}�9�8��u�f��j4?�E(�������|NK���b�z'2��Al�Ŀ�j����5~�o��C�Y�+B�n�R�8�Ϯ0�g��J{�P�h��A�.gHs:���K��[��y�����g�И�L�vF�����#��C����˨���Dk��v�nm_J�	��ƕ�J�����W���f�A!�3�3���brk�����	edS��ǯ]���6DR��e�y�����gZf��~�F���ti�e,��9lF�O��O��J�mXL~�㋮��!1�ά��ʖv���#��zP���V1�v��
ٳ�$*�2)ˑ�q�����ۆ	+�H	��p�	%� w�*��Uͪ�����'���ػZ���"�����PxU����5�^�+ ��?%~��+Dg�3Y����sf�����m�G��	)����k0폛G����0���8��e�T��O��`���Fa{ޛ�ov�1��Bׄo����\K�b��?ҥ���K�Y*!��]Ze�^�����Wf�V��l�o�z��N�Q� ���xo6�oj��ΐJ4t\oB�'2h����dIj�:�c.kg7%wK:t3�@�@��W��'w����RS�z��	�_G��B�{�+[�k�0��VA���M�s@�V�#��Yۮ!:}{	 +t?�0߄e;4�sߦ�L��Q�'�]��f��멛��#����^������f e�N�4w�C�	;����#L_��>@�ց�R�<YФ(�߃�Wj�W�:/��o!��1-%$�Ŧ��
�д7�h�Dof����"��R,�kk�B�񥬩���)�tb�	V���[�+�۝�8����և��;�`c"߇��V��-�e �&��5V�>WhB	ha��mZ<�Y�띚��3��<V�����X����ܕt�>W�C�` ]���0i��(���|!/<�)�p3�UO�md���a����Bo����؃(bo�MD]�@^Д�㞰=����80�d�2A:Ӌ��|�zs*Z��r=s�_Xl��I�'$V�t�qX@M��:�P �D&��&�����߀J��]�Xpb̓T��L��n�da���Qo��2[Gf�mM��Y�M^�$��y`��*���;`��ޚRLǘ7���:��Y��9e��
�3��8�-҉E��A{�6#}H��R�s4}_"ξ�>�:�a����?i��!J����S�N��4����}*&�#���љ-�|�l�7VzJ�u��@(�-�Ge�Č�T�>�/Xa������y7m���
����y/7*�"�EÏ�����Y����rl�4H<p(;2��킭Il�/��잖6�>i��J���`���!C`�S�TS��-y*��Cb�\Q���nmdL �whU#��w�^>��" o�!~�@~ �y�e��	n�%��]�8��/G[�+�C��ޕE����ԟ`28q������D��iY	cR�H�I��ݗ�X̿�)����]��L$��l]��Λ�#�q�	�3��^�����:J	N.S������o�	O��п.'0�C�]������u��U���#�_G:��~)��O}�[A"���P���6����̣|��0=4����$��%	�|�M���5�R��.�9���W�J��c�L�ӓ�eRs3>�H�15$ή���^��7�;��}� ����+��t��ẍIw�Ȧ*���-��BS������84�{#Qu3�[v��MI�=�@@#� 
X����-Ϋ$]��E��7�g��������pd
�V꒛R�¿���E��	��~�'������MPn�1��/�I�bB_�El��]�u2VYk1�B�	@5�x�Y�Y}q��?z��'�KA�[i�/>>�V���Tzj��ⴞ%����b���z/�Xz,���]�븯�yzH�D���<���N2�`4A	vQ�'��1I�2�}�s����m�,p���/�	��Їw�y�ِ'�s������``Z\����DK��w'��_^�X+���+XJt���5���+�s��/��@�}.�����;�#�0����=\f�T�7�X��7U����M"x[�p��r_^����8f�|�Pa��Q9�q�{k*�@�������QH[kl-�f Ծ����W�s`+ z!4?�6�5Xlg�[�yz��mZP��r��lߓzl<х��Vkm!��,(E:X�Q����&m�n��X�Ϩ)�˱(:}K
Ηk�_�r��,��'�(�;���(�N�t8p���H�E<��ߌ��=ڝ��p�	�Խ�Vc��A>Vo�)�3�l>�$�qH-�զ�2�k��$.�M0�1���ߕu�\�D?��m�g����"� �ߕ���Y�	 �y�d�_���;�{Mv\չ}~$�"�I���*�;�@���.��k�b#S��ׂnX8��0t���� �q�z�,9떈����刣Ǐ$�]��W�����.#��0��xP��c���_Hc�*aE�b@<���<:-W1y60�:�f�l8Z�*���O�4�{�� 픦
�r��gr"�k�U�*
n��>����7�)��iw�����pfmU[7����ZF�EH�?��k����h��J��U�6�:�J�zX�i���!ȝ��U!k;���&P��G���p��������X��<5��=��'�?jO}��6|r8�M�
�՚�����׌>�s�t��nE=�O.�!����9f��(�=��a��`���uWRg$"�X��q�x�r�����̛������p^
 �c�&�)̘�2�
��#|2��ge�Et��-L0�=�ʩ�æ�b�����Е.;�V��xM��$u#$RJ��,�_���ڂ���#�ĉQ{w�a��H{�3��h�!������9OEYa|��b��~U?�C�u�3����ˇdHS0$��#��9�����X�i���
���FF����#�s!榥��ٳ�(�-Գ���v�2��r|8�N�S�6v�жr��t�9��L4o���꡹HMi����"�!"��.�c\�P�z�r��(%��l���� xpm����D��oZO�[R��B�)"2�i�e�(�jK'�ڧ��sh�IO�Č�]5}��)���dn6_�G70�_#�*6���9��{�w�1�0�ׯ �P�_8R�����P��K�+c��5���}jpA��<C3#/�C��-L��B��{m"ݜ`s��|V��W�C���&��i.NmP���� � z�/�˘s46�)����e˪��z]��篥sm�[p��4�2���]X�ӭ��1��J�F)˞>[Lȯ���S��+��
� ?n�Ͻ	85�«$0ϓ�i�
������ ߵMeCO򜰈*A� =�0<�īs̜C_����9����.*u���w�&Ӿ!he��>g�̏���fcV2��%g�	�RK/�������N;��bd(�@ei���X�gW��(��ɇ�o����u2�逑��f,3l��i6�M5���H�-�	�.u
ܝ#����v�e�r�%)[����l:%�]���}�[���G����e���8}C��=�t<���b���Q|�[;����T�d�~�� �E=H�(4h:;��w&q�+&��\��7��j�O2��1N�L�}>q1���M�µ���h�B���*���P��~�0EH��`��k�%�	{�0(V�[@.\��j�xс�e�vz���<m!��^^~�.�>4�xwg[^�#�l��5�ި�6�Q[N[�5�Kr��߃�f{m���]c��?��T���)3��C#a������!WPN/���)��M�aE�/e#y*����I[�\V��z&�%��-e��+]fP�y�y�\yy�/(�4{'��$���"����G��?ޮ�䟲��$�ZM�#׉p�6�T)���x�<�B_P~g�D ��D���Ę�`˓Ĩe��J��K��@�l_�c+���p���� T������yB#C���yhj�!(����
~~M���ͅ8H���~���h(�P̏z�jU$���p�z�%k�C�c�}��\�;�y=�tx�ȦO��S�4-�?��h���O��1�ȩ����88t�s�?���4��0n��D�}5�-$:$q��P�HTS�9jtI�i>�R;�Ī�	�>�[��"�vi8�e�K{o�Q�қY0啈|��3dS:�dRp(cK}iE�����h��}�c��`2�h`�y�J�t���=���F�F`�ro��Vr����m���J�%v�BVX��I��_��@W�� ס�����IM�;?r؂�j�R{4������Z����%)@�cbQ��Eg��5G>{0p�_��$w�qb��L4�1�Sp�m��2�1�˃�2s��_�]��:os�(���*�5��R�4�#�T/k�5���`eD���A�)�<#����*i� �8%)M+<�)�v��F�
RE�����;6�dn<����� 0����lҌ���0�ٳ��~o�q��k[���9�񎁞����޾�EҵنO{J����H1�p�G����P	N	f7Vdrm�#bk�Hh�Ӷ�"ԭ�d�9�!�c(�-K�XI!���l� �mkf�B����.��ۦ�qlI-;M�R||���ldLsT�㙞/U���@M.Է��]��B`K���D��Ev�S'U7�����C[��+3(��i��z�B�H6��
~fb���.�Bc(���ےc�1�şn�UR��K��D|[:��� �"CO0 �	���,�4��5G�I�l2H���.�ϟb�Bd��������}�L�F��㻢FI��y(���4�z I�	e足�L꺙b�x-�����p�a=0�����I9���pJn��g<��~X��;d<Β41f�c��S��'��&4ľj,��R�1&�����y�R���`�W0���\�)�3um�'1�$����F���5�Y��z���h��ַ�3�ПBqE�0%RT	*��6�,��;r*�C�� ��b�Q}���Cˮ�b�Ȫ��{��~�Z����-��w�0�s	�M�Q��-���vWҍ�-):tW`�V�0K`�xB�dMT9\6�Q���z�*��t�#J�Hv�$O[ 3��.)���A˼��D\��f��!���nK�*���,ϑH?y ��@�'1_��3� � /V���#+�n��V&��J}����=s.7j���K1�9��������g�37O)=q�W�����DA)s��h}��w/{a�=>ݨy�=�-�\Ʉ%}ʹI5(:�`Z;5M� �Ɉk1<�z��kFZ��N��.�3��--������G���}zR+�:��x�jpS��X%��G����rw�w}�z�#�'�pU���f%M�����fk�&1`�D+'�ɩ-0a~q�Wd�EҀLC4:w�lBo��)��H�u��_$) R��S���_�g��>k̕�+�̖ѫ�x��T{?�FC ��g���������	�<L�.�Y��c����RT9b�q�F2��M�S.���1N�Ȣ�JNE�������I�<�F;�$��A�_����oᜃ�|�����a�8k�>���~�B��J��*Ea*i�ӥ��sUݨC���Nu��Z!+�I����]���~�`&�8�Yݐ��c_ �)����8���_S����-�&������S��hja^� hTa����Ծ��;��r�5�~=�^��ԕ��V,�&0'�o����EI���v��z.����1�=7/����������u���#�f�����b���i&`wTSb�X�)��4J�'� Q�;�Y�G��x��fc�f�(,�6W�	���a���Yu�"+�����<me]��U��o>ν!fO%��H9r�"'&�z5W�!	�i�B]J|.��ׇL�<;IȔ��Y���H P$�LNykM��VCnn�cs�ū/�λ�^H?W�,��^��O�/�pa�EE
�Vː����A��1�=Xk�n��HGL+�.���-����ZAj���NA�=p@�	�P��� (U)bu�mH���Q3������̡%lj��h�"��ϩb�ʈs������UHCRc�P��=w��w��
����ʻ��9��Ķh����]��9��D�C�,�G�=z��9$s�l��,�z1o�-Q�jV����
NJ���/B�Xe
n]��IxI��=6���G���e-�na��=ȣ��^���l-�,�&�Im�3�-��d0��o��RЯw�r��x��%ݯ��{��E�k;�f�?��H���J㜋�w�ڀR���L�`�B����ge��.Z��B��_��Fe�+X�%��$��9��<	T���+�%N$����B�o^7���kB�M���Lu�K���ms��쭄?���Ϝ�ߟ����O��TtGG��a�-E��s��i/��Yr�w�\�͖�8�Gy"ϛ3�����p�e[���i�-#��\pc
�F����GnMi�\P �4&,-�c�'��OZ)~y�QpT� ����Rx��@�o5��,Mo�߆�?7�b�"�Nd)
NP������^��������i	H@�

��]Ȝ�vV����&�(�p���x*I�x����v�f����p�ǜ�n��=( ��N��OL��I�ݘ�E-b���珙�X?n"�/D�d�F�e1��p�:�=S�n��Yk��'��=	�$�(���vkT�Q��'���˱��Cc���K��!vc�(��8�3�73j0�m���F��P�%�<�G�j "��W�K����9`�c��Ѳޒ3�#�K���l1�Mh[ȷ�Z�M���7��3Z$�tdӂ5d��ޜr#�����6�G��>D��-����.m�5߻��0��.&�����&���\��7U��)"I=N�6i! CD���g�l�\���2ze%���^lq�U53%� J�$�T�%�D��j-E�&�DM8�xV��42��^Y���R��u�p�Z$���L�n���'�h#Ŝz������M�$����� ¿��uQ�o&H��"k�h̢�Tj�Q��j�����vm^�oˠ���̀i)��7jw�u0Ɲe���]2�R,�%\�E<N_l�D���6R6���<p�,�!��"<}
fVr����T���X�&	d�f����ɚ��U����>�+�)�^^wǭ1(᫈9)3~�$w����]�:��y	����IM+���P�^6�����&��O���70���t�L�S�����P�OM����i��Rr鏵���j��H2l�\����<`�*
}p�d�qP���T����,����u@_?�� �"q����7xm}��-�<t2�����۶d���O �+�v
�P�6c��@N��"0��n�e.��Il.��C���G@�֒��������QX���h�����s�Y��2�<����ƒF�����r��q�����v{Y��&X��y���ImA�aN���U�'�$�h@8cP	�۩��>,p�u�6��c�W���"�Gz�YA�Jv|F�C��B�¾%�g�+��u�:��V�
�E	,
B�E�;f/5uP�������~�mML�\1��i�%s�%~n�@^׬���k�d ��ѣ���_j�`@�0,��1��.����YW��DO.�	��a���ʚOl��'�̤�bM�K�����l¦P��b��^͈�W��� ��=@t��Jy9��,]#��-����5+d; �bU�`��l��
�[�_�4S�`�Ъ�4��d��7Qz�x��F���Zl%����C">���g�LbJ�iY�W�(D�6f�+tݟ��W*v��7��9q��<�6:�|�_�T\��zIv��|J�7tZe�^���D����-�q[�Ύ�o2�FF跌E��� ��Ukt��`�R{���.�[P�C���}�t�m�X<�!myDċ
f��p�&%ʛN!)��,i��	��X�
��-��Kސ�0b%)5�J�ú�們�d9�iKL�,\��r� D�Dt�ȕ��q�3��.qg���&���8���>�'2�KS���uh�ٟ��<�q{��LΆ�32A�1L�߉��+.���ӂIR�V�+x�/8���j�p�BUe���&k�D�I�%�����R7�a�D�B	�������Bo��HD��WH��S�؂T7���'�<.gRQ���7����/g�"�h'p��Y}9!��ERH��[�~MSl��ϴ榬��_kc�b��������+A>ڭ&W���i]ڌ���k�6�N������ش�-+��s�"������7�&O���ls}���WdIA��̕�f#Tt�#�p[(y�<�.�_R��'��d,v[>�P<r��o���QB���Ά|��0lx�[�1�q�UpJ��͔��y��	R|�T�מT0�ĿY)�X^��VK^T~z��FV�H���[��!U��}:��-J����Y���-&sKe
U/w!�J�����H`wà��&_q�E�WU.C��W������8� @k�RӺ���F�=c�MG�Y�O����v�^���<j*˰��O@xn��oPW�?@�A��u�?�ǀ�<�Y;��Z(���S�c���_����9��ġ�U*�V�C�'��2)�De���!ձV-Sj?�����Ɣ�3ӷ��],f2���P��L`�?�%�
]��v@�6���ۦ��V�S��������u�P:r@��)`w�?Jd�QQ7��߬^���-'/R���XrN�xj�f��*JG�֯��s��<u��)Ĥ�'���x��T�WjԜ���k(�T~��!�ފ������8���|o��{ы7&��mHa3��} K0�p�3;k��C�#�I�4�-Ũ� �]�)�)����OL�?[\���MA�'�@TH�(���)���L�y� �u�����K���y�ד(�|��sƋ�΢��?�*�D��!�0�tTdp�ﾩ�h�I�ɲ`.��Q�N@���/3�\���B.?��e�N�!S5��"����?HQ[��h�p�램�0����rYc�9B���������!(�o� -jJ��1i~�͕	W�6����1����u�įD+�	/��&�_�H��1'��I��sn�O�=����،(־d��Ǖ�C�*�^mw3[`)޷��,�sɖ}A��{�6���c/�I��ilZ>?Ok`~�|�!^�0tWn��s�1fVmNkcݒv�u��<â"K�V`����Y�C񫤱A�ߣ���ʪl4�(-Ef�ٶ�&��OL�����;��զw���-l�R�XT[h�	m5�(d/���0
1������p�eQ������P�X�ᦡ��C���ޣ�ì���ua.�#t��'�U��V�y$ɛ�E�b��U�Q}��b(���$b�u
�Tոy�dQ�~jc�t��8��t�IG�R�
�W�-� V�=�3� r�v�x�ح��}������Y!����Hz'�#���]�ӌN�D"�P/v���6۟�fR�`�T|��sfQ����5���6��hߐ��nJ�Z�
��{;��q�ջl�����6�^�Y#y�3+�xje5�*u��ާbf�*m%9�����Р���E�-�J"ɼ��"����f$���j���'���t�EN=�l�a�FR��7�&�2�v���R;bZ�zD�,/Z�0�:~Z�����d�I��!���F��+��v+�����nG���6yFQ|�� ��
Ԁ��+�y/2�rVX�[�8<���֭g�g�k�x�.��;h���8w?̺O��U�c�"���0~����1߁��.�Qړ�ߣ��Z��~'%2[Z�W*5|�u�����*A��>N`�|�����Q�'}���^�مc�����%�/��m~�U~��i���I�f�%ˡ��FɁUkjn>�b���Y[��?��9
wĚ�A�o,��W�K��a��ѕ*;��^G�
*+;�*�)F�Ѱ���Y�e�]~��'��P𪅬�����T�V���O�yd���v.M��_LB_�\*��[Sy�{vZ��9���_.���$��r�
�xA�ƃ1�4X	ix�1l�&�tg&�?�xD�Q"O�RVN���xsp��js����'��V�l�[�����_]%8D�I:��Cq[N�=3-�4����Ё�Ƞ<�4X<j��3qkW 7�!���4o�\xM�l#����9�lY�d�#R������U�y��N|e�L�g���n ��2av��x��YP:f�6�;�m\�����b�^�'��.	27�Ix��m~ɩ�D��aC��L;{�{eԗ��nAU�čH�t��-BiH]��z6JC�����eAX�5 6d�񳅧p=��R��Ք�� �	בW��A�_��upy��'�-.�j<�-�]%Ȧzs �~X�/�>�?4�Ak)�QLm���X&ᶞ��\��<!���b�c<G���*ND�����hc�&z�N�;���p����������)���ul�q�^����B�GmowE�!3�@���7�b�t��mrn���"MdZq��Z��T����l�KO~���{ڸR��|��W^n�#ή�г�s2m�@\�;M｡�����W0��(ρ�T[���	r�>�t��b��\�)
�w�Z±
KI�1��2S�a)���w��v�1��X<@罘*F��[ؚ�F-�<�����XA�q���Q���0r��mP����M��HZn���%g���b�����V�F���&�~�`\��Rz7��8A�^��ׄim���C�6~1�g=����T��;R��r���{X���I}��'����;Ժ�A�C��jZ~w�F���ZR����;�Bw�t�3�!R����3SjM�KX�3���Y�IC�I��03���r��5L=yj�^u>)��'�h���ġ�S�+�� �jwE�ό�Py�-�D�ec�K`��K��c6�	o�Rk9(�GV�7��&Ge�Әa]]W�~0�k��v� Z䓜�\x��<B$\l�}'��k�����B��Ǧ�#�ZT���8������s�0�0�m��
F-u>/�[���ϕ�RH�g|���c$��Tq�D1� ��w�wq��DČ�@�_9��6~�s8�����>���p����60�4�Q�bm���˫7�;{�0����K�r�6��7Yj}kayag��:5�ZV�K>���3f���`��F]%�Ta������ݻ� MaL	����fdl/�4Cc�`�Y**�_�چ��p�O��{
����Ic�/�Lα}��>������7�&�V)��sm�8�F��x��/ݓ=#H�~�{��d���d��n7��dqþ�ޣ���h�=<���|���t���'͙ެ�5�:�c��X	�.%zf�[�,�}@��.�����6ӗ���Ϗxn�C�G�~av#.S�����#��ຣ�}�Ր��6q�_�M�E�R#&h�A��T�F���,�U�L���ֿ'`#{u�t��f)�~.��C'���8ُҌ�_���-�/"T��;�o�~�K�$3[,�	��.s��<���X;Z*rz�LOV6;�LFM�ml��b7rS\��z���I���#i�|t�J-�e�8�Ř~�WCyY?��ㅉ������ʎΕPU��>@��l4��,�c ̩��2�)�8%k�(��d�=p2�GP��U��%�%L�-���G��^E�&��
@ "������sB��þ���g����s������F�s7��K"x�D�HL�;���I���^�& ��X�!:�i�VRD�'
����p��"R����^P��\������g$Ʒޫhv� p>24b�\8�I�)!�c^�N�	�tr9�~��Lf�b��v*z�e��;a+*�uU7�y�M�.k��Q߹���ď,��%]��18*=Ԉ��?�_ǩ����w]�S�Q(�B�w�E*��I}��x�-F���\���tYS}�"�Bڭd�}I#��w]Il�:��JR���b	�}����ѝ�t;9��t�D!� j=K��vrc����Y���̜����.^�)�]ʬid�GMY�%º%���ʜC^�����|C��!C�W��Y�9�VY��wuq
]�l=��\�Q�t�v�f��8��+K��hI������.��������LO�a���[K�y�ޛ~��Ǹq���պ����蔰a�෹�L������6���YW���ď�Tc�wG�u\�fq�N�ָ��5Vw�7���(�&YPo�ܕ��s���X1��ǬgZ���l�
�ĝ��>���,�9V�iQ��(i�a��ӱד��d�����C�j�sZ��U�p<��@ �O��j�v�vVV��|��6�(�	&d����D��f9d�TA�`8��WK�f�-(K���be�?U��A�;Zn ��F¸&�Ъ�����w�%:������ѱ��W@��J������T]����(@��-C�-�����6$х^�^��i�,3cy�:g��H�31�'�8�o��QV*c�D�P��ta�L�vCf�]<�}o묛0�����T��+�
�E��4��ܻ\4ah�~-�㓴�������j�$Z+`�2I�+*��R�TQ֘���6���A�9V�Ƿ>O~`�y����6
�aܱ.��V�sW��`;cΜ]gi���O"��,�x&���t#�.�F�f0��Es;ઍ�4I��ZH�X�Z��`��G�X<P�vTV�8�@�{�;�S�t��Boy_ƯIbq��;m�9�ut�4�fB�M�1&����Mpr���9J��MY�fC����ݣ�d��4�yt�k�L-΄[��.��D��yHtZ���S���I$(�֣w��1��*�:�D�F8��'ĂзOw١�u�B�����J�u�0�8�.�t���o��x��\q�7�a��kKb2����U�O���l�x|_ҷV����,TB'b��2N�"�y ��smw�ks��כ'�΅a|����v�YH4�	jά�UP;����A���31����
!$ֵ9���#+�g��C�>6!����%�4b�����0N��������k�)Z��\�l�NL���ɂ@SZ��w%�"9wNx0A_��SZ�N�;��#h�y�0��6�y��$ѻw8�%���	�C�R���_t3�U$D(Za��(	�N��W�����y�����s�·3�����tӅ��}���C����R(�@���}�%�O	�R��lP�jd�%IG�)�f�/R�)�g!�����_D� ����5]��n����Y�b�Hh)�2�d���?t�JH��9�F׶�������@5�;�͔RT�c_�3���Zϊ�9��`Q	�;��{L#,�Q8��,��#�}aNb�ΒZ�S��T���� ��3+�i�V�2%��������zwQg|����������ȎϽ����s2z����8G���[$�����so���^d��.J�;%Ԍt����)i���sm�a��`�h.>v�!�'�ꕫsBztc��p��E���E�hX��7���߀7�;S݌����a*�S�ʎ�Jt˱��&�ޮ
���&����(Ѝ*9j��-1��Nl~<�0�u8ji����,�^���@WA?�j8��4g>d�	�8�`3��?h�/�9��W����}gW����¶[�@���*�F~y	�Q3R���r�{N�aK%�ܣ{�lC)�={�gQ�a��� 2JH���`A��5㞫d&��I�3l�R�76w��M=�J��U�T��
<�(

ߥ�࿀�H寞o@�/ݦ	_��j��g�Lj8���ݜ:$�u�>��Y���������sk]����x.UK"Bċp��qgeH&���f�
�%�%�Ȳ.Nq!I�1\���	�ȕT�S�t��E�����}�*�Ox(��:��_Uj�ݣf�V�Y�I��E�&sx�I<$�����+9��F-�	�P>���/�Dw��,��3Ǌ�?�t���/��7���s�����3�-�ѣ�f�U!,�J��^������V�#*j���n�*���o"�tSk��	���6��[\�����8~kNϹ��������u�\�ƪ���}#S�f:ǆ�3s��{�>����ZD��v�#(�l�`�?��
�~1�O�tS�S#`���`�
��?4�Ma�l9��@γ�g����7�r3�y)	��g2� t^�c0�D��'D"������\lʅ��_kLx�����;?
�a	���9g!�� ��5��ʕ�\��$y��nF�h�/u�D��׊:�]l6ә{�Y6�xZ�Mb��M}�ح5	%^�x��(�����1�[�5Scs�-�
������1�dh�|Cxq��IP�&~�'-.[�S�VVE7����^$���P͇�-�ZB9���n��ؒ�0����!j~�g}��ܬ[���i�`ʁk)�WN7U��u6�"�s���"��_e�8�)�0Ɖ�0:��zT��Ï�P��R��� #���G\��E��'��-�z�kω]`�A>(��+���5W� ǣf����+��ŝk��^�T�7^��d�#LYf>j��`�cxk?�7B]���AJ�SY�ʰ�g�-/�[��(��&��>0胴��r[���U`,��:�Ok���6A 1w��]��9�4V{�^I0F�&���^�5�)P��O�p�y��@�5T�ٳ~�Qjm���_��I��Ny0��-�ߜ���#�ԃ1�KH�j�0M��73T��j<�J�
kM	�\��<ě��L�V;7R���_m|3S�o�w�f�+�kᰭʷ��B��J��2��������wn������y�b�g��Z~Wr�B6����i�G��>kX�lލ�b�H����{���}T��+"+��a�+�Y�O@ύ)�� ����~^��+2�(К��M��m�m������G�}x�5�
�5�0s���O��q�P>FiG)F���!v/J�t)��5�>q��.3���MZ�\sV�
��"���|�6鰄�&O�L�P�_AN�W4.���K2!n,���	+�n'��D}Ԯ7JQ������hYK�������1E����~޽��۸���+XK���\��Z���a�8/v�Kq�������Bj|�&r�7ڨ�q���E͂\��4����9yɫ�@fg�a��o�
%++�N�}�E6k�aX蕮k��j���~��Wy��	�C/R�п�8�d�pA+������:� �R$��t�3���sp񨂊�g��S>������Fq�b!���k�3������R��B���ɻ�r+�9\��x۹�������
������4;ݥĒ4mc�dz��d�݁ ����q�R��M�I��P�s�«���,��ES��S.��mvL�7�:!q��sx�=+Y|�~��O����.��ʕ�J@.tf+�I�N�..�A��e�0�Q,H=�Cf�M5�K�7�w�p�%�{�5�TG�@�F�Wm�bd�O�/�"�J�q+���K	�M��"��15�*�k�������W�n~���zC-��Ԕ�An��/"ŘmE�
�?��Bh� ����}%T\�A��Q�i��	v"�� q�!������:�O{z(4�=�g�m����p>�d�-��N}g�H�i�� `N����A8�j��N�&|�m\%.�KBN=ԍ> [_��%%omh�IY����b��_���4��A�juc�����5�z�>��PD��`7ә"=	ʾI�P%(W�x{#
�i�lm4�I�2��Ym��a���SG�����U�!ֳ��	�)�*j�7�6���
�tP�h�ڸ�i	�"�Xh�:��ܻ�UGv�Ō_�9�5�e����I�=Ȉp�eP�����Q�����xwlN���\��
P/����SF6��F�f����v����
� >-I�4�3��=; l�CbZvk����,C���@W��ط��k#��o\��/?n�ǲ�:�J�����˟L��K�j����+F%�f�-g�[L��*�����<�;̎�W��p�d>��Ѐ:`�
����6K�̒�}A�gZ��ͻ��̘��y��u^�ET)^M��w'� ��Z*9�rp{�[��>��~��a��ќ{{K�7���	�����d���w�"(7��Ҟ¾/.i��	;j��ƈ���|����������l�=�`��mv�}��O�&+4�����]��H�U��v�������M�h��L�XL���3
vۻ �R���W�����r�&������ߗ�M&m�9�P0���;����F+HO�>��E_G��$��{���)zrx�΋���94~��q��V�_��Gv�b��aS����a�T�0R6��(\Q��9R�T�/ڗ�4sFgy���v�^Z��2V��bLb��Q�L�������x�5Dűֹn����Yf��������AJ��3��V��n��}sH�F�����A��(S�΍,�Iv�t-�P�+�� |�����}�rte&�n����Ed��
9L?���h�I���f��u-�n����t00����^$m�1`i�(����"�-�̒^To/�������U�d�sT���� |����-����μ�9?d]?�R�7���g�<�����XE�P�"Eh����$�Y5c]E�+վ�}SM����V�o�l2s>�;M5ɶ`{؍�#U��N�4�����f��{��n����KW���U��$�h���9锤�gj#�2�s��Y��`s�f�40���Uo�m�('�)r}������j�����t�u�gy�ks��dg1�N@�Q�~�⨾z���g�i�l8�^H�h<O�0�>[�=��f*W0���]����x�bī�.]��8��7+��R�v�ROB�m�/�G�N��s���p���B�j��_^��p�|�l7{���:����)3^�3�`��z�Ia�r�\�������5����sYJ؛�𾳘�W�3U���T��K��InY����f�oɹ�:#s\p���C&]QY�C�i���t��z�&�Ŷ�?�-/�K{ O��P���'.��ˀ�[\ ����Ss:e1>eW�0L%��Y^��Q�OTI��֚��"�aK����U�#��A�kn�����	���z�z�+&j�n^^�m��T��<�3�B�Y�.۷����)�
�M/���4�37, 0�Hj�����l��Q�f�#az� zՄ��X���·���s�7?�fs<W ^14���A���A,�����B��_NL�/�F҄=�Q��� �=DBO
���fE=�&��W�?T��`_�g̿�w�3��W*�Y��d�X��Ew�ڷ�Q~y�����Zba6��	�l�N���;�#Hk������`X*t��U�+p)펭�e�� q��X���H���.�ꍷ���n.�>���$�q<��q��\�SleW!}e�d��PD���'>#D�D��A�aަ�槃�,�Kރ,n�u�M��ʬ��{��u��p�S�<-�����&�1���G��`B���Zt��f'G�%��<#��(���_l��&�ҥ�iBe�`�׆����0������g�q�
���H�#qN#��K[D>������ceK<R*5cr�U��rhKr���@�_wb�l�=�KX��^6Nĥ����5�5|���CJn2,���!�t�o.\�)\kt�@���8��|�9�驴�M�6�"5����^-�� �}H��I��!�։��_~���8�]j���g�����S�81��z�P������F�#���p4G��[*�4�O��8=���--'v�r���Uj��l�}�!�͸�k��df	��7קt9���7|��p3��Ѐą���I�=�\WSV1���ΛQ~^���o�^L��6�.��H}k�^��b���{_n��)p 48GR�OxC�Ҏ6��"���0ǻLl87S�5��aw�\B�9��T��`��u�OE���r��ɳt0#�Q"���չ$�K�ј1�r.�R�w�>���p�]pM-YO��oAD��?1��O	��[n��\w�*������ҹ7���caz{�7�y��A��"��e���A����(��vU�� �I	_a ���T��~���_4��T%@�:�_�0 Mt�ß�P�i�f��o�Ǐ�h���3����]�)�����~��,�Z!j!�]Q�/���ҳ!WpIw��xG.̿�и�'��|����|�����P�[죦3������NfRǖȽ+�2Q����;�P]P�l�h)���·0Y,�<��ЍD���^�.���&����ؽ��[X����h��h������Q��,*��-\K0!Tʿ46�5��pˣ� ���&�Ґ���e���-�[^��%���/;,�`���+�l:$�1����,Fep� �>��Z,��=��;�,�F�
���/|��s����!�]�]#l��?��F���G[��1V/B��dy�<��P��4�.lO�Qw�m��s	�M����Q�0a^]����˃\���WB�k��\��F�="J?��f޺Wf����x0KZ���À����f���R{<8 �U�z{R���"_-�9<?V��Z�/|Ͱ��SXDqCʶ�W����a�������[M)2 �)��-q�vrC`]x)Y���<��6AKJij�/�Y���#аN}��׊� 'Ǆ����/njA�JH_���]��+v��g*��5����,����$N�k3��e�n�Y)u?~���2��W�g<�vH�`_�ߍ7*ր����Ҝ�`7j�M,�N 7���"�*����D��i�ʦ��".%�	8�x��!�|�rO:X����?�)L���"�KZ����oO@��l�ˀ��a#*yX�T7g��%��B�L(�;���O���K����;AEyX]Ɂ`�#��b(SwI��h�����l��O����͐z7e���œ�q
�Y�q��B�vX�ZLk8(?��b�X^~T$]X�+5�3��Bbҫ�
)T����˕C$�7�Gޮ���=xh����j�J(��� �`�d{�<0:p,X)�bA��&�>��Q�&����2h
YAܜblݺnBSqլ�
�t�~Q1|d���e�'E!�%:�����Ď��M�FZ\��.Շ?�/�|R�kn��z;��$�,�ĺ��@Y�qB�P�ȎT����N�a�ʢW���K򭃤�W4[��^@�рT��B�#�A���6yq�C�.�,C�ϖ0.(�9P�CLi���������[;�f� �q�jU�5��N��[{�} t�׉Hgkg��L��n.TXn3/�����o|�T[��!c��N9$N�z�P6Z-���?�m�Y��*���Э��GW�ڌ��w����AA����5�kh�*�����E�|�e�Ӝ$��w{�� IC\���Y~j\��1
�"�TB�&�p�ǌ����U��[���X��d�o~��PF��"���X���ܳ�F9��`J��Y��x��Xƥ�/��nK�r+Zt)U�c@_F(;;�fc�c�`��^w|���w6�����kEߔ�W�M�� ��	�:A�)��Q����im��,� ����Կ�p�nu �c��T,�Ne����W#���K�1�g�D���ڥ��"8D�O?<��1�����v�T�X%���'� ��2/k\��L��}���m�e�uRR#h���@��,x�#.���ޢJG�̑��u�]�4@	�6���u����Č3ˮ�y=Z.I7��{�\��b<2.0r\3�s޼��H,�@dD_��9]&@�x=�S�jZ���A ��!_ c��[E��0����kb���с�oJw�"�nR���s�ݐ22���Lq�l<��*�BW�y���� C�l/��M	���7���P\���>��Z��%��>���Լ��^�u D���
��&��'��Zx'CpQ����O����_H��p��?��B.��^�,��>�|x5˟�R�^��*@�RT��cP��*mFX��4F1\��,U�bI���W���f#��@�w��n���#?#=~_��$����y4�m�: ASOp.6k�R/lف��;��ri��B[��|�����UNU.J�S�H��KϦټu��L;�L�x�s�_k	%���I5��Vu��>�bb�=���W~RS��.���R_��S)	�t1-��t+}|3 ؞�Pcja�C�'�V�2n��q쫸	�7c�yb���T�Ț���Lɾ�KB⅝����퐐������b�V0�m
�3e�]A���f�$ۂ�����T��,1�������we�}R��+��a�u���1�%ɖ�G���T�c0a�<(�����*�Fd��.&,랶-���'_��t�]��̌%*q}��~N��4�U���uգWK�2��t@�b���
!Q�gN+�`{f�/�/�P���{_^ʩ]�e�r�%%��
"���Jd���^�1l�a�n1d��8�`�r~tދ�na��>���]��ş 0B7�gd^�W8ING�DLV��w^�d+*�~5�Gr���/��3Z m>�1��Ó��p�&�P��(�rZ��u��
�� ԰�_NSe��TCMr��>03�%y��p������ǅ��h��o�����S3,�~��)�@ھ=�#@��Z��I!�X\ǟ<��@�������Jq1ÿ�CEc�C+���l|�3R(fSFsSo)���R�',9z.�{�n�\ئ��F�%�ǛvUH�G��N�^�\^K/���ԝYCNۘ,��U!S	,�[L�7��$����ke�9��6�D�4��C���V�,��P���ց�*R�����6��/2���㐄���k�����Jz�R{H�S��%���c��?�i����\����N7:hS(�42�U��YZ�x�J���RPוGI����"�t�K,�m�p%MO����P��B�T�[8X1˲AR�|b�Fo\�H�?�P%�5;��|"��{^�[­��{�W�6۟���*�*��Ֆܚ]a����c �*]���v�
����)7<)</��������`��kF�|IM��E��e�>P�{���փ��?ڜG6���`������dӫ�^�'X����U�G�1���C-K��،�գ45nĵ{���MÐ��� 	��`?�̨Z�ӐD�Cw�,�$]�c�6��7�[�B�K�P�D�BQR,(�Z�;(��;I����0�6|�1�8_���T{1��h"F
ؽ��˺��}-�hx;���Y�@ȱ�:�\�����;�ƍtso>d��p\(+5m@m���������Ӗ��S��a��+8qt���k
nW@��Yre��]��F���X��#hl�W��y��8X����*�"Q�D���z�ٟ0���=��T�$��{x'K��Y_���u ݪ��������20���j��ZjʀPW-�Xg��A�1,Omك�"�XF�m`���5�T3T6<��2�g:]�f�&�C�ڟB�%�B��������<�X�'[���?8���W�
T��:�oIPy#g�^���d�s�E�5�Q���Г�c�M +
��-
�iCl�?ǀ/|��[2T~L�a�2Z�eǞ^ Mi�DPϰqi�芍�V�Xo��-�ȶw��Ŵ(��)��YeQ�iL��on۞�G��t��j"�ShXT�����zW��?��V���戚�$�-�;�f��7�I��������t�����x��X��Х�t�tg�=��Iыay���p��Qy��t���v���Q_���n;5��b����
|m�r!,^L��պ/�~"�����H��C'��O�nT�f��oe�?�@U�����9"H�p�x	���b���)ˇ���
]�H��T'���F��БD%�6���ّ��8���ͽ�$ �e�����of�(���	���T
\py����[����o���7�X�wW �18���+��%��a�J�q�a�8���I��#��w
K���G�$��8��u���16��>�dbVuSk��m�����`�>h��;ۓ���o�Ί]�������ۼ�q���#/�&_:d�V�9�VԠ?Ad��;�g-� �>ڨ.g��W��k��504�Ƌ����'��[�:�F�bX�oQ��tE��3v���,�
�ͩ�:��b�4�М,6��RA��J!:�z����j�5�7$��P ���'��Nx�p���_hٽ������&N��r߾��`|��9���0����\7g5�ьm�{��kt�v��/�3�UMa�Zo���|żGVx��v��c���g �'K�p��ӳ/��to��yF�~��n�(X3b8�s����Ux��؁�c^�J��L�
�H�
��l��H���F�xL�E,�8n�w�m�t�*�s���<6��J�+��@�/����wB�~���D���S���x
�yo���eNQ�I���f��L��Щ�����P��������J����̕t<	K��t/ZW�t�<I����3[@�;�H/����7��Ÿ��8�\��=ƍ�PK���K��_�ݠQ�hJ:z�a���$��`L��3�&@��D����lx8�x2�:�0��F"n��
���L׫�A��V%�?)Zr�P��t�ȳ=��6�ל;p���Ј�p���N�N�����j[i�k�������\�y�ůMsf=�]�ag���3���67m*{jw��qk� �=��(J�I}��+�2���$骩\�G�`e�
hN��5�$��H�f�Qf���DQk"��2.����v�-�$�92�oC0<r�`���rV98���5wc��U�}tߔ�7f���{ҖXZIa�$'E!)�9��\[J�4����ic	�
r��P@�����`��}����]J����1m��^8����/v�vj/�L�W�LZM��}*�WT`������*�7�g�p�` �.j��dya�؞K�7s0��cǁ p����4���z$������4k�;=����0�(��S�M�<m��J]2�iЫhjki�ԫ=�/-������tgrc�X�B\l����ʠI���������%$�3�	��5V9uUU�-�[��n����srj�4{�F�fco���ɦ鹀L����"=��b��XU��$�y��6���T��ғ��F��Zc:�q�xI�v�o9��� X�i|��wr{U����P��w��Z���8{�k�|�����
W;��Si�	l��z��@�9�e�;�ӝL؁]Dz&�'��g��/G�t��4c�ݓ�����$�DF��uڛ�˼L$0N���rӨ�^�>����Di���ӹ�6�yVl��&�抳�����B�@�����׵�$�9C<{ĖִRF\���\և����B�WƦsР���Pt˩Z�J4�(�yd>���/&X-�Kz�5��6���%>������������Q��3[��=Ѝ�~i�.zle!�l��l����s��;�'S�ĕ*I�i���-א�?�V��;�����%���4,�*Ã�z�_^�I��5������ȷo�(|pce�F����.���͸�*9���-�Nee� �q¦]�+��w@�(�J�/�.I������M����͊԰d (͑a��[�U��]mK��_��r�It��>M>��8A�_@��x�,[����������!z�t�_��]ŕ��d[�[�*U#0}�c��;i�Y�PC<�B��!�`SKlmt��*��m$���ႚ���ԩQR�r�8ߠ�yJ��o�m��J�<���Q�N���9�2J����N~�����"D�䙱�R��
��U���[��.t�!�sj$i�3�}@ܗڂ��v&"�Y~�`������>R�D%ǚ15�7�f��Oc$��+�NP$��]��+G��Ґٓ�bϳi�������#�e����Sqvzy��bc(�\�Q�(O�]����ˁ�����I���e���=���M���5��g��"f��޴Ʈfp�
TD�<Y�&����G�W� �pr:���fI���� �C�˾��:w��ّk����� ���;ҝo 8�.��0˙y� :Yչ��H�l�ُ8�Ŧ��kU [��V��	HŒ����\�>��Y�6�g��8̦��Za��>�#�x(=��a���75T�����g� �#A|܋0օ ���_¦
u:�z5�+�um�	�n��݄�O�dR��t0�Rƌh�Ac��V� ˅�zE�.M��P;xj��u�Tl���F�������uII�֟p�⟗���gi��_��g��Z�ন(��%\�3<a"oX�T`��?'�{�+�+�t� ��>�y3,�%��m�BR�݄-�㹉�e�g�N��`�`A�T�FoM��(�Y$�$��vL�S�,��?LQca�l��(,%�Dڅ&�z�@-D�}�"��2AG�&b�Ź��o�\���F�8!	q�2��Ǧ&@2KV��4�����\r��R�����\�����8(�x鼑��?�Ig4T��1KX�c�B�P7[k��=���{�˳�'��o�E�s�5Y?O0R�u��۷'f��vU�6��s���\�޼�H(�����E�hHɎ��@��R�~:i<]�/�]����*��\+E�E��d��.���P/���k�5��:�݄-��e���b$�j�I˓���q���"�F1��Y GG�ӨX�	��=.[������?��]U5�.���\;6�8��w���RC�B���k'��Ng$	!�[�p�}P2��@ɯoy���g .Ol�@x��v1�[W����RIJ�W�L��]R�ށz���i�ݧ>L��`q�!{����H���m�XTH]s���k�!�u�3_$O�ݘCF�|rf@Pfì|"��
n
�h�	mՐlu���I��"x���eA�N�FF�Ez��`�"�9�8ډ��oB�[���A�o+�[^�zC �.)N���c��âPӨ��h6!-�A'�)ݷ����W�W��Z�}S�Ʌ��h�z��
��_�8���W��v�I����Q<|eV�V������(���+����%��SD	��Y�[���%I��5>���on� p\sv�D���<݌i-�7Tx�=��U��ă�i��n\�u��XMabD�RS��T��C�z '��)L��%Bw���Lz���k�����f��R��Kb�����צ.fmMZ5LC�)�гH�d�*�H�aq�K���v#�#-�U���xV⏈sP$�?�!%;�)�o��CBL��E���|g:���9�|�EN@�`D��3��O�	��771���=�Q������[-����Qn6��"�EΚ��{V�CN�G?`A\�̖�̜M����ۖ;�b���i������E��'�����s���R�;�i�p��P��.�o�'qr�
!&T�[���`v�cf���*�ڐ��I��2rs�"�6a��������I�$�����b�_%&6~LHR�ƙ*P5q�����#:��b�V���_�_���&&(��ս��ir-�N j��X��g�)����K.��
��:�-��bɞ#g��_�����sZnԧⓄC�Yl��K��뀞5Uh��s,�es�5� �`Vܝ��!N�i���WH�yֶ��$�4a�.1X�k�6��v~�(i#In��i�>��e�3�
O�r���C�m͍�7SsI^�z_@0Ƿ���kv��-X�C5����+o�hv�v�nb8n��.�L&����G�%#���غY8���P?�n�E��(y�APK��+c�
y��x8��	��9�|M�ӑm���I�C�H�m��+P �Q;�S~����?Þ�,7�)YS?50--�3�@��t�t��;�}�.�����UVc��;���?1|��s�5�*����
m�$Tؔm� �e����.|s8Ǿ*(��w�ˆ:m&���kL�5���A�m�6�Q�{)O�8ߒ�F�J�h���r�;ۅ��/=X;Ͷ����GC�^H�W��{��p�!�u��� v����m���.g��$�R���)�ZI�u�,5S:g�0zJO��FJ�X�f�0ႉ��O\?�l_�ٓ���{���f�uU�,�`�J�%h�|%�=�2���IfH
Z�~���˰���y'�Ut#¢��4G��Mw~Y����>���v���-��4J���b�ѢuΏ!�N$�@Ӭ5{���vJ�����=�ŰM�Jp�Ňw��K2���OX)�r`(K�F�
.��DJ:t�_
SE:��U�1ʜ�W�q��yۺZ
�Iw$��PS*?�W��2��JM�0�}��Q���\��6���D?+k[�Gn=�"�O�c1�-<6_|'�`�"B'|˙�{���C�ӮQ��4�h̯��q��!X����c�oN��F������{����W� M/�3>=��0:B�mHU���ۗT�P�{e@��F�P7�����d& �p�g#'ь�Zy�g�@����ڎ��lm�16��h]��֍�ټ�����c�Z���rGS-� �����X?��!�*_$������~OfM�{�zlG���B+�˔�~B]�r���iAqzΥZ=�����T���}�ʏ��i�y�BX���|X�9Q�6�ٱ�

�8�΀��":�**;S�"���[��!�)��a�e�m���{@�#�m7w�2/5�f���m���%s~�[�J����A������R�f�1��DGd:��N�읕V�0e�v��s��&>!��:�\ip; _��v6EX����lƦ�}[�G����O�e>�0�]c�׽��m�μ�P�vH{C�ǭkF��p�.q'-�R���������InW��_E��s��K����t�G�+�"c�</��Ÿ��������k���	R�V�d��A	��vZ1婿o���!�^��Ʋ�'>L�/[U�)]�� �,R����c`�cf,6����W�Y5��׃���h�>�sp<�QQ��V�:3~2h4 T�~m�kemO���AG�!Բ_�W�%{K`�B�@D�;�ǘ�����.Z�h��M��=�)�f�8��۰x��vِx���ɭ��yr�]��{x^"Ԣb�h�X�M�vwR��.w��^��C;G���h��*Z3����Ŀ$TT�O2IW�U^+�T�Aq�kSf�����7��ԧ���[���С�H�1�32�Z=��J�Ė5�\���!Y;�p�
�mT@���:aY��YT?4$E{��NI�W�c]��ӣ�c�'���_����N|}�Z��몽�Z�}��bg3��������]L��D
��O=�P���;���bx�#�J�JEA|_:z�� �ш�Je�l�J���E�3��m[@�X����dl�?�����:�U���8˃�@����
�^������O�V�FCy��o�y�9�8\�އ�F��buJK�~e��z����%b��{�+H%�̈u��W�J0�&�٨�^�eh&�3��/;�G|*�,����E<�'�[��J��U����\1�רl��oS�N}��g��m�o���si.��)��089Y��Ql����:�4D-2��x��4=d��i}h65��hȧy�g�y�f���� �Znh[A���m�����Nr0��'����ߨ	�'ϫV���1�C������M�,ʂ��ש���]ȋ����>�z�������p �T�.�#�� �K��� ���(h�	꺍��z�JTI���V;����1���y�K1_�@;�[�b��L�zv��WBN:�<?�g��t��s����S�Fcɶɂ��<����\�����I^�T�B|��М̥�h��'�ܟT���^0�)�RoJr�`���D��e.��&f���\M��< �Y�g��u�����EP��k�F!���8�<Wr��3B�*xP� \��	S��u[�X�Y�A/����
�מy�z�8�0�V��+LW�*(��{�0E�>�eE�J�L�ߣ��&�pl9qU� �{�ތ�D���F�����b���p[�h'���A*�f��Dd�������č���Ɠy>�`���/8��K����S$�ī�Å��]�*ZF}<7n��6�8�2�Z�`�����6����T��o��΂O��v�R��F�V��w�@�~}E�W�9S^�҈���-^��%���s#a���F�<���&}�� b%�]H�q��� ���ڏ�fTx_�o�#'Y�Ӳ�9ڿ`�8KǺGO��J��I�!L!Y&�ad�-�6)�p
����s��"�@�3D�C ��c~zz��&��=��Z6�*�|�q7U�r����8;_݂~��G�p���8k!��j�_��0��O��{��oe�g�Jv�j�Kfs�J��C�s<h�^�V�tO�}����eh׏ 
7��9&�Հ���8�����+��[8(y܈ѓl�˫M���roR����6{'$x�`�zI\>�&I�A�?2�[�I^��Wjb��q�(Zfq�z���/���-ͩ��L&�Z�?y<a���@$F<���G�
�%	�g�����E�98�~���x.�3�S�R�qNݳ�ǳnHZ]�����6ĺ\Q(�v{��*^K`���ɖ"��_�� �.��#1n���%�W2�"_�/m���!/��(���8���A�W��r7��!��� ���D�
-�S�ʥqF_�����ۮ�#
'��L(�C�Ej`�x�Ջ�y��-����HS���� ����M�g4o�	�)Q]�;���p�=�q��+�R1�l�����$�9:h"#9�4�5��h'��J��5U׮y]���=9���*�t,g���	�@b��Q�~�PC�V�4�pV�����RV��ڔ��~u�_�m�8����`y5]nL7�
�{�{��r??��	�cA"�	i،�	�@�~$w�~��Y���)��3��P��Q8`���1�A�.?�S/�f�f��e�+]h�u��&���t�����H)������w����Ս�^�Cm�Ց6�EE�jŃ�̀��`�-�%=Ǉ&�f��Eq�X���9�s�{�����N��j�^�V@g����g�^�m9Mf�~��a���`΢��<�[��8���]Vj����<Sߖ-�Rt�^�另&lD�#0A�5P�̀~6R���l,)���|���/s���}�m�P�J�g��`�6�,C�E%���b��N]��2Q�F�Mb�J/IFq ��1�v�mB�����+���n̅Z�'��ZOrXc]I��2���-?���1b�J]Q�Ѭ{� �cuy������H-�>���t�=Hh�|\���\�r�^7��J쇈��w%3�!P�u��4.�K �GS�R��F]��v�����!����ڃ�� b���e��_E���\��I�
������p��߾t�Yե��A��Q�Mɶ�	�&=�4�������f��)�G�9J�B�3T�6�Shm��ocU�	-�����E�WR��<�m<IR�$ S�g��&����F�i�{���y��F��9��w}��L�����7�yǔ!V�6�o�c����K�g��2�t��Ah5kaD��YŃh~s�q }#��=�9I��l��ߟA�v"s:Cɥ��TA��k5��A��w
�s�9|
?7��[�g)M���s�/��; �y�J6����^��6���)���{-o����xUU�<�� ��R��%��'�c��IZBi�'v���9��z��%.v�� �ǃ�5����+�\��R��!U9�Ϳ�`Z�X� hJdŨ�Jy�*����aխ�W������"}��;�|�n����8.
���Q��s���&[o���� [$��i�re�v��H��^W�����R[F{!��-E��ރ� W6��NgT�8'M�m`�{��=9�G���"�1�*R��-�:���s�/�>}�����OY�irS��-2���8�.���!�1m&<������.#�=߰p��eCr
ydiTi�=�kX��F����*��Ǹ�hF��A����:
g8�ە�T��Y�rNs7�Zk�8E'���՛l��?5Z@�Ҧ-�j�7��_���nO��R��_���DMB�UikY����-r���9Eb�E_�9`�N�bO��Y����B���.|T��%舘, ܹ��3�i�ƨ�#��~	�(歴ZX�L킚� �F��QA$ٺ�@��x��<6܆�E(�b�؍�O��df@K]��1� �A�d��+�#aȾn	���VTIW�X_�w����{6�^`R�o>�Gt2�Za���тo�B�s| ��Gr 8���B�N@{F�P�C{r�s�����c�:"��'�嬧Cb����qa�E;_z�X��G���N$��g%�4[�� ��d3�:nN���8{��^^�2�E<���c�!� ��CSL�}�M=�c]2"T�?���"-�b�),�Z]=<�yN�z�v!;6�o���?�����"��i����4!���`�&*�T���/3��0Z4v���\``3������f]N��@No�]���ߎ�_z!���_�V�r�bZ�+
�J9���X���!J
!d�]�:���}�����KR�_t��u46����"�D�q���A_����/����Ҩj��a�.���B��π�xwm���i= p"���	ǣj5����<ᨼu�p7a	��M�p��~p��q]Kk������`�����!ǯ/�jÂ!u ���Ԇp�$a����<��F�z%)m� ok;�VH� Az0��bhyy��7�EY�
ݸzT��m ?�L�	����7���JcРE`DbU��¤J��������N[�F��RL���P��9�eB��Z�2���JDT���
�(^��.���DEm#����q�&&�-����&�C���г� ��f�UF&*.=��
Ze��=�R��l�4-b�.Dr��w2ކ�@��z��!(W�x�Ktka`j��X��zU��2&��*�j߬B�Fh�s;�iV|tW%���;tC�]�h��R��y���s���I�d $�V��w�{x��&h����8��}�л�+,���)_��f�"	42CLMaϐ�%��3�a�N?'��ޯ�`@���@���_7u/ ��&�sW =�֪�y���j�tő���H;-�"kV�Ć)M�ё�#`����0�͝1r�|M0��9�_�.��F�4U`����Z��S��ږ$�X]����P��
�N��By$R�Gjn�@nF��E�ٹl��Q�)��!�����9"�NՄ]�ΚNdq��� �ƥ��V#aRk��0&�?rU�NI��ܿ���;]*����b�;�#&�3!�)Q�����,����!ͮ�Bg���Q�a^�c�"�2(@���<<�}�r.o�FgCp��S�^5,�(��b�1��IKEX�j��dϫ��?*��qv3/|����f�%���1;�u���|A�Q窝.6J�h�<u�u��_^�O�l�	�Omþ��>����A��?��2�4������`���E̘��е/uŨ��Ȃ�Q��S�&|`�Үq_��Ҙ7I8�Z?�`�S6'��8�J@(��Lfy��s{aR��&7)SN&�v`�^�-�2.����~�F��5�%Ϲ����E�굇}suȂ'�BҞIP�ܸ����O����;�^��U�ۢ�����͞d����v�<���t�`��Tw�}�!�(Bk@����f���|� ek�Z�bc]��8lj������fG\Xe����c7�q?oN�r�eY� �<s�q��8D����P�(�ovf7��{Ab&L��`��w�w^tM:@��f'Ph��WAk�����[;�}
��Zy�?�%������R*��mu��L�l �B�/(��d�g��z��͡��	~P�>0)Wձ�o�G-���%�sOx2(Jl�:��ĮbN�X>�F�`�;���?�����"��m�P3~�?�-�W1��?��UK�5"�/���^ ��h��!I���ܷ�&R��nX9���[��f;�{�m�3̬Ov��G5��W��ɮ���RMJ��[�+2}�?���{�w9���3��yϕ�|�� �b�l;Q��s��<��X�XLTɆ�'2���!P���v���]���*^��|�m��hӃ^G/�*gB(�  O)*�t��R�L�겻�޿Y�Ɠ�Ŀ���Ԋf׶ �X]�z�{@[һ��E՜NzC���� K�(A&�M��1}���P�'�*����}���A�q�鵷�_�l�̓:��A��,	���/���RC4��p{kǸ�1UG�����QM�s\���O��j&.2��E���KJM�:À�2�q��U�s�����i�防(���G���ɕ&�BP�~�����`�3�p|�����7���R�2��J���� FOJ4��컑m���m{���P�u2[)~y!�-/(?G([��4�?}{������GyF~'u/���%Q*�Ga���@E߂�OV��H�HLj�n�m.r�RS'���,�|
���W\.�^	�2Oa>��2B|�3#�/L@r�� ���O��T�=�b>݅��g����aO�=���P�$�h���k�I.UMγ�!�ﲾ�SX�5�!�C�t�0ʮe�߲h�z�ٞ�fv��㶣�����-�w��Ь�X����E�Gs���-��z�ݜ5���N�r���1��`kkU����NJ��T�Sm ��q�~i\v+C�S��v���u4��߹T�ۗ3��Q�H=���}��s�+N�{h_"&�o��5��Qvۏ���^��e~�E]��G�^L�J�X�N�ddHw������/�.*�>gK�ܥ޺H�긻fR|�Έ��<�>nթ��ٷ����6]N����_�_�(G��)a��_7"m!N��Z*�a^��ƱMT�O)��3,�k�8ͳ7��?�"�7�N�<�:�j��bn��\�%V�9tWQ��X;�"\�w������ǎ�̜e���w��y�㞙���V� G�,HWs6�fS	wbe.~�r�y�c��\�ҳ�b/�o�����lx?;��?�Q���̶#���y�����Kq6a���q�_���]�����(��&����"7O�����'ǂ��U���0���0���v��6^	S㰡J1�]���V����j{��;�r�>B�Ls�����-���u��}5�
\s.u-^�ϻf�K������y��+�΁�})y���Žv�̅�y�������*��j�t��*{^�ӧj)V�ɩ�؎y�[X�%��a~FRn��&�Ƃ�L��AQv�S��R��L�⫔F�B����6c�F��~e���}���|�+e�S�-gF�T��$f߿�w���	�x\�:��!����0?��z��S��S��y�4��5u��uL�ɳ�9�Gǥ�L%���[������D�9]�ԝ���1"Q����|r����u�"i������%S��M;�K)�	���}�>�9�,[������iۀ/|i�iǠˍ�(�e���e1;i��t��H��P@]r0ec�M霍�,�V֙��9[G0n3�R�k���z�ӛJe�ʯ����j�%"&���T4�� ����ɶ[�4r�,�r�A��R��T�.��"��ٻ����8|<�< X#;�vt�O4���(�}\�
+{}���>g������ʅ�W��X�T���&Q�A1��=/�şȤ����}ꯜ]��B�9���=�'_ǋ�@��8�����)&$ʹ�&�`�Ao��=�W�4��!`{RGSV�B"�OP���د�xϛ��1=��C	�η�jA��|K/W+�;@K�r��:ּ�f%>C�R'��('ͭ9z��ςH�
ja쇍�h#�o�4'E����q��Źf���?���mL�^IZ	�{�Ag��$G[�s�+Qj|?�r�sJ��Q�	�P$�G�N^	�����e |`�@�w5��������2{�B�Ls��}3��|c�QsNq�_��|j��wr��^DO ���(d�<}]�!��_��O���2�����J<�q�zؘR�KZ�1-/%G6��C����f�!�}��6k��A+dxGJ�����Y���Tq��F�d���*[�g�����^�M��8U�����f�5�K��XGY��� Խ{%��1�p1���Ņ�,��y���/Ud�!,�$�Ҟ��s`�h�~�F�S�E���F�����x:��|��D@�4t�\~z C�	;�����%�р��`��X����:���^O����Uz��|glĘKp�zg0���g��"la$E{O�{ᩪ��M��ٖ`�^���&�1R���-�g�i�����s���ʝ@�S)�]c�-�WP���Y��t�p�3Qz-��a�����P�}��ԙB��2�L����dr��ȕ��W/o�����h��� ���9Wh�Ag���iN+�[x,�Tl��+%"��D߂�<�L&��O�V�[/n�+|8\��А���Kb��CJF7>����E*Ԑ�����e����������g#�J��(T��A@c!Mp��!7�����c��G�O�� ����W�3���r��ac'H�beQ8m����%a<_�3�$�W�����e�&)����gT7�#��G�&5�L�mG���g�G&1��u>1�P�Y�\�V��[��SਁWbΝ���桓�x�NJ����N���y$�q��=)Г�g�ɟ-�=���ew�5#�Ԋ�4�e2o$���_8�:�3d�Wc@�p_/3��w4�k�S<R��8�W��\붯�k�Mܗ��t�Ӈ�<l�0H��L�jS���b [ʪ�d�Q���"�� ��h��0����į6`�}q�
�h+���*W�8�����Cg�&��>�k�?�B<4)*�݅�E�ʭ�XՔώr./����S�D2T�3������U(`����5����t�+�z��pI�N�1jXч[!�>Hy	2�/ �3D�W.����̈́j@j�Ɛ�3��l��ʞ��f����E�b��J*mTR�o$���M<��{3P��6���k�7K0f���d�K����>��!����`E�������1�t(���W@��l65$�%	*���ُcj�����1@q9�s=�K?�*U������d1�~*�Z��1�����?T.�����<��K���'
W��g�W��:�r���,
�m��M>"������[H�����j7n����ʐ���>�@�q��[>����N�f�fW$S��oqi! �
�l���!��'�Չ�cz�j[��X�B������V��V��}�H�f�D��)"�����Ư��-u� ����Gr�/��
G�)�qY�5�0�T�K�0��f�=RgUwQ����S<pm��v =�%>ڇ�l�d�E��S��W�/(G�u>��$�Ous���5<��}xd��l��y���J�&������K���%�⣸?YE���O���^�rdl�]9^w���PT���`����g�EpT�U�G}֐)��-1t(kBz�о:���ؕ2^kM����)o08y�����`f%��\�D�#�a/�)���D{����i'����W�e/U���R�;!���wT��6��a'���  G�\܌&��u���,��	������v�.It_}M؛&�x{He�\d�h�JdӠ 8�)u�|vs�q/�_�,�~[A��I�1�H�2�����%o#@�=$�&�ρ�n#?9F�+�)�9N����He��1���6����t�=5���gˌ��P ��aa�ʞ���l�.��E^���L��% �9���M�Օ@��~~��KPZ�� w߿� Є�<��U�[�z`R��3����c���4��h�#�����8�6�Ԗ���2��aJ=b�8�Ӑ���۞�[X	A%`���6@Nθ��UB/�T_�Q	��D��xPlh�Z�`��m~ c�N���%�w��l���1B�k�9j��f]i(�K1�)������<��N�fQdӏ�L������9?�hKs�߲��a���~��g2}�$�3��LB�ܛ8R��A��UN}x��鍌X(�XlPz���;���D��M��Wk�1?wf$��ErU]jެ���^.f�b܊`��q�F��X�SX���w�� �~���ı�]�e�^p��#�����������d����O�/�K�g�	Jۥ��i e���J~f�:���t�اW�fDBY�6X�d3�����
��"�\B�
�x���A�����KDU��� ;��
�V�}c��K��`�4�[������k|�ɉ	?� ��l���@�5�H�����摥%��)�n�>���׹kC�)��}"�������������O�����7عAQ�]�ʅڼ�	rNba>�Ҧ _5z<I�/�p=�flp�_��	Bޙ`Ļ����#�а�!��s��BA��Y�6�Z��2J�޺iL1�N ab4"}��Q8(,��&{Z	��2�����]v��%G�J��'Q���ԇ�ۯT�3�R(��{K��H�|a4��ZՈ���K\�P6e�{(�ut��]��.�!;�F����٦�P��5X!��m3�1Ѥi#_��f5,�6����>�!t���^F��)mX��hϰ���T�@�&�;?H���b�7')�1��nP��<�:��~�������Y��Hn6��v0��J�!�ה�o����E��U ���[�����ն��l�Cg���=]���~v�Yh����
�'��a�[gݗ(�*(�yv>������g��5^m�$r)��ȃ��Ř�BG%�N��0���0i���b[%��%(Stj�#0�Բ�w=u�iVK�r��q������3u�>Ѓј	$�]A&q� 9�MW��a��D�@�[s{R�6L鑶�Q����'$����}_E�]�CS�"�$�jw���K�t��Z�e��\�!�(N�B�2��vu�>0G����cf*�JJ��(�����_�yI��߳��7���g�኿ G�#m���c<���sW�Pd!|�A��Q�h�v��dYr\g�����Kp�e�H�R �x[.�;�(^,�A�g&� ����8Y�V1>�}�>�XdU�qۅG+�y���~�ԋ�[�'R��rE�q(i�F�Z�6�"�X�Y�.����n%�k�q���A�rDU������;��J��	���6<����Z�D�N18|���e�����G��vÒ�h��z��.���3Y�b����Qپj�]%���3�T��S�$�(n��w��,޽����ϸ�"n�B�����A�CF�<�m/�E���W	����r�N�0KUj%�۵�H�	w-/�\(~�%_bUP.�{ݤ�J2Sn+�}e�T�bs0�j�j��5>[k\{��֟ۀ���ް\[|�[z�3a��ٙ$�;���~��{H�o��#�ϐP��Ī0��q��޿n�u'h앱��`ĴK.G��T��S[�����*ʺ-�n��PƐkue+�Z+m��������W[���?���W>(�:�T�&�1굿��Gax�MImx�l�'�E�&`���8r��^G�a�9���.��ͮ�U�a��4��UP﹐����!_�y����IT_�Fet5&3f��KYR4۰h#�x�@�,�e mNj�?��K0�s-��wo�>S������HX��>`�c�h���V�Z:� dǃ4�|*+>�;�j��A�8���%Cя�Q�r���U����?/��7��/��ΧdD2��mF�R������2)�󟓅x�a/��jLlp�dVL@��1l��M�`ؐ�*K^,��*�v������Z�[��P&�VQ"2�$�?3��e%z���̔�2����c��q��䥟x���(���6��ų�\� ��a����_5�R��'�e>�]��ן�`}߉�R��+p';� M5��.�5�	��qFWX�X$����*4 su��&��� �F��=ΚӰCS�_���AN��g���Q�N
E�|5�`�K��Q�8�p���w�y���qe '-zw5��✽����Y��[

ۅQ����N=���׏0?�I�f��9Ry���ê+o9G³	��{��ϖ���{O�H�����5ԥ��"���v���U��(;�ҁ7h:�^Y0��]�x��㮀����Mj�Xκ�%�����7]��~u5ܕ�˰��ݰ�&eP�������Ը���`
�sz4 ��G�vA�d
m��� �x��`)e��Di�1Q�w�v#�5���g��G3w������"r+��7gɴ _�x^��䭋���5�b5f��!��&��տ�mf�@�󺉠�:&@�
A}�/��0�_��c�mꗘ6�F��w��(�=�n����m)
��X!(x���Q"M嶲#��Sm=���
!���2��c�B���9�w�z#n�&���`5?㡍(a��u����	,��Rȑh|4'lo���zo��N���E&�T���M�q�RTͧ��!��D�@~Ұ6j��@�1[�K''�]?�ܫ>9����E
?L�D4'��d_��"sO䶃���c���4�f�'	#�}�ZPށb�r��tHkY�Z$_E���1 ����F�@����bݔ$-h�;3�� `FD`R��U�>� /5X��;	�zۄf��F�=�-m�0���� ��8i���ٜ{|����J�>������w��?����d��z�Y�	�L�F�V�Fj0�c�3קnL5�h�}�?[3���-J�$̦_(�������P]_�Ec23���{�#��4�B:��lCu��*��蘩?:8iw|�G#�5�MP������FS��܊HɅ�-��QJn�O�{"T�+����~ǔqW�dc,ˀ|�T�u��=���E���3�m4��M+5.���
-�"�η[��i�!���Xi�k��Y�q���DL���'Ltg��Z~ujh���ڭ�_]�!q�ҺZ�p��m1����8��i��� �iE�cH�&��{��~�X���l~�+�l�b�ܽ)Ӻ�<Td+���Ĥ��4/�_�oێ�+�_x��S]�z=kG4J����B�7����zY���Snȷ�����_�s��8�0�����'õI��C��%&T5����_3+:�9������W�i��T�R�ү��Ҩ�]!��y���,��3�j�E-���W�1в�U�b탧#+��O�ZC�C%��}*�y�?�l~CN��z��(�[�l�����bŪ�HO�iFD�\TE�	��^�->��n�ބ��q�����9/����V׿/n� �T��F���H���a��~|/W�kX�6[�Y�d4�)�M^p�P��	��x���7�Zȅr�z�^\n��Z��B1O޷�@l�^�ul�d�rQ.�R��>#�rܕv�~�����ҕ�=�ã+�U�D%�
���C��%~M�CPG�i�~�E������k~e�\�ȭ[9�Ñ=]��
�Y��hfr'���˝$D �u�Nв����C�e%����=�"��L�~����68�Q�S?2��y�<~���W%���(ot�]�ތCX1���%g���&㴆iڮ��ݓ��Z~���컒ET{*Eh�UN�3�剫ߞE/B�౪7�nz��O:���X��/U�Ʊ/�f��3�|�6�=i�ᠶ�:�x_�E���ԪHNd"8/u�]~��ܥ�u〠��6Ix� d�r��|6�� &��|�un��� �r���x���l���Q)��pZza0rP6a�H(tE��*��<�UV����Ƨ�h�kS���Vy�by���������Pp<8��G7_M֙�~Ӧ�͑�+ٹ*�}�Tn[��-��$�)�r�=-x� �]��ƽ��6��Z����c�k��;�eޞ6@-7Z��
�[�\X��+�_���R���D��"�0o�{���OrX���� l--X^$m��>N���!�e�1du ��(Ic�̗q��OI���wND�/EN4����#x�W{%��E包Ԇ�3s�ĵa�Vn�����q,��XA��� �>�7�4B"���+�x�1�DE2%i&~"�&�����g+>���4�d��`z�RƜ�z~���Љ��zQ����da�ץ�/E2;�0`�����b���?�b�O�$�34����F��H��Yr��P�Z�pכ����*�����f�Ŵ����dZ����.h�S�~�D�I�$��Ep9M	R>X��5�^/�}wF�¼v�Th���ӻ<W+9�p�byǍi��RA��c�כuB�1��`�K�)k�gV-8x	�c����i�EIv�ñ��@���s%Y$-������P�)��R���=y@����=�D|t��ޔ.��'�	*��±x�e-G7ʕ�� ?j͇¦�w)RI��ʺ`�ԢZ���c��������Ӭ�v{�A�D̝$�wz�A�ivC=;@���y��l?��=1�֮J��M	)����� G�?kҔ�TwBC�����w�L��f��Q�H��Q������5�\��5�ȕ�x�ؾb{4�@�!�Br�����r�/=���tt [����vO3��4�|P��ߐ�]�e�Eў�������q�7y�����b8��t�ߝwO?aW ��^�t|Kq��t�H��tm4nvY̡��V��9Sx}{����~�:*��L����[��®�A���O�yT���2ދJ9ޝ���P���>ܐ��V��3Ty�v_X��K���Ro?��܏�[�S"�v���y����3A_�1D�%�����FR�K�*�O�h`����ڔ&s��\M�dQ��hD��X���\d���l.�����.�h��T�'e�֪e����f4�ęK$�2cD��/����u�l~�N�-�y�un��\�"�kr�*P�cfpz���J�F�:fQ���������롮���U�jo�B�i�[
�����2��}�n�(���K�g'���"T�DR��tt�1����n��9rnV�@��p)�(9
���{���:���0L��j=c��iy�w�.:	�ejm�7����=�8����e
Ԅ]�N�AI
�ed�f0n]��Z4"Ba.қ��a����!�#�6Yh��#�z��Wg����>��/;����+���*�D5����؃�t�ׄ�T*����c�V8dL�|*�D/u��dw(#h8��M��0V@x䃓n~%m?���#©�v�>
Ⱥ�2	�8���%���e�����,-9���c��[�8`L�R�?�b�6�b�~��K���3�&8�x��s�<�w�ج�G��X�C8�2�����/^��z�ձXbvSF�U:�jN=QF��E��c&���#j��n�J|t�뇭���9(�񁔤@�rSSX�U����M��,�P�0�@�����b@d�Ï�Z��Kl̚F=M�Ѐ�9Ϟ�O��q�N�߹OU|��?���#���<OA���p�`����=6�����#�U"��]���b )6*_�n��6@y�)�"�;}�I�&2�t٭���u/�\'g,�7#�?�&��u��&gFj(�d������U_`EN�?v�b��r��;E�[^�K�ClIy�'鯙�=�{Q��Pq
 �Q���$V�XƩ�H%��Ktس��3�Nl4�3f�*4� ���&??	�+j��V(���\�f����2�W�g�^O�5g��a��Z�m!�a�C8_YC-�� Y1LŬx��_u�5*w�D�YmK�rfV��1WiVLY,L�ံ��E��A���KGC��m�{����s�_���n�HD���>p�<�0�7�����K׭���A���36�BIC�ẻ���৩��uG��"z�m5!�:&���*�)�j�Jh�P'����5߆3�L�~n�����{m�Y�@����c(4�]փ\�8��/�¶�_��<��󸊖t��[��d��d �BA彨h�<̇>Y*��׬S�/�Y����u��q�� ���b|J����f�{f|��;s0s �b�Ƅ_��b3)Y9g鞂�-Q\������ʆ>�[GT�<�'���S<����f�������Jn
�#��_@��u����w�1��9�t_��[���8��R�$Ǣ��N�Q�P0��|@��Cn��$׀���A��tBN���f�5�c��������;���e��:���t��GѬ~�'&�0n��Υea��F����g��߽�@EW�D�X��Yv�xk������۠�<��u*?eW��"�7��7�
�-zI4�:���U�9H��|�P��\��\��7.���uZ/�x��҂b��_j�8_�����V����|��נ',�;d��i�ץ��l<�^��ȒQ�.D�@Sc��k��1�U*6K���
"�)�h���밤s�/�1ƽ�j�q��N��UטC�랍�b���,�X�m2��6w��#�*N�f�誜���@3��0�s�O����Qf|S�S;%�!��%Mz�2�m�Mu��c���oo�Es';�qӣ��D�EH�$��7"y&�������v��:�T_�E��
�}���wcE�޻cЅAe�ܭC��j���?e J��E`#47|/�O�I;H��Yo�0�zh�{t,m= _�S��{��RH&Sx1k��b�q# �!��B�I�fO��H��Q��م���Rh����L0BЫ�yO�y��퇋,��?6֝����!�q�X��a��Љ�ct��ʁ����&����qE�A�Ȼ�O!���Zj�ܒ�=%��)n��l˾<dD��5i`� ���#{�W+�>ّ'��o�n	��v�mD����4B9M'�/+s��p�EY�Rh
���w�~w��g�o�9G���4�'|�������^�:�2����B�G�Y"y���J��W�jr�O�R���������V�x����؆iC��#����V)z���}���*���^�rm�8L�;b� �����;�o���c��J6S���.WQ��#�f�����,��JO�lwXݦ�д{7�`1�l��	��揇k9a��7�!0�"����Ƙt��֓���\�G�v�8�}��s��^�p�tj��ٳ'��I���ŒwS�S�銢��j�=�cF0ꦈ|'�\z$���daQ�� X��0���<-lR!
+��޹�^��"c� ��QUn���#9t�9�R\?��Ĉ�!�z��(��.���;��LV'O圁����4�U�PbÈ�?Ģ=�=#�
��ޔ�Eߗ�Q�i��tS���+{����{U��=�T�C;[f_�z�,r���[`�~>��e��{��È������=�����]�JF�up�	s�<�eZs}2_��Fu��oq��(��Γ�N��,_Z,h3���IU�}��1�)�-.XP4��O=������8�rf�5�Ou��4���O���1F����~�����4��O����_Z7�d���/�����׸���I\��,:��9�=��a�J栱X��ęɅ��v��C��io������@q��=�"QQnY2��qV!x(QL��V"���Ԩ�oz��
�9����4�,Vl���p��bu��k������0^�=2��m�*:�뗐����,T�l�g�{nt����� 3ـ�k��R�sV���4�ܺ)mUW��qQ�Nl$�N�Pk��ޮ�9���m�ub
�
��v�@�_rOv���
A-��]���]���!�b�8{����2�\g� %A�Y�?VxJl�D�ss9���`er�<\����<�|~�,����F��f���͇a*�Mp��:�Ъɻ!"�X����#.����z�Z=��L�A̘��p;gx%3��MD�A��
����%�x�9�	N>o{��C�$D|���HN^L��ܬ�4�(��	�ʯ�,��/J��s�>��B�X�X�#`�5�0ψiRW��NŖu��D�*7к�6���f����Sٲ�1kP�2�����\�ms��*Z��+G����O�Z�x0�)4�q��V�Quf����D�I�3Ⱦ��)Kd]�ɹ�#��,	�}�2V�Z
���z�]Y�6~_�oք��:�$�汏6k�U܋��x�r ����� �1�o[��VG�к���"� �=����u��0h �=�nUa#me�+��y��QFob��S��bF���p�?��̽�%Ӭ�EU�g����3�\�A!2H���f6��N����@����M|��|r(���/��h���2�e	b����G����Ԝ;�B�����p���q��v0� � ��>�$vGH�9��	G�/&����JME�b��%ř��W�K��Cd8�5m6��]��k�?;��-�bج�K�YXhTc�9!���\�j��ڹ���a�R��P�}����;�X1x��c~� ����|OL��_F�x��m�r7O��wt�+�`�K�sPPo�����.ejB����<=�����4-�C����Hx�K��ƀ�GS�F�,l��6�`�ܯ����z�O!���J�}ƌK��κ���)쾖��։��蹕���1
7F�G�&�͂�(O�f`;LN�<��_�J?6�J�.�h��Ų�2���F�����0�r׸�}�~���#7Rf�P�|�6�|�_�8�����CF*]c�|]ہP��V@Bl��#f����J����.�Iy?F����懖�h�돺f�[&3�;c�R�ޭE�;x3a@��,H���'��Z	\Nj�;z�� t�_����º����<��N(#����Oi�
���64���E"�<.��i�+����I��k��}qj,��� ��'/����[���6����5 =BfaJVk�C�m�$��Eizt�eSM��R�qUL���z`�,4�tX
��ꑐ�b�Ruw�%"M�Eu�h��G8k�@�:!�?�c&f���ٔ��]�H��=(C��=�\�a#�Ì��|���g�ͰS�����H��G,��4b��6E�a3Ca�o�l�af]Zf.��%�R� )��~����Y��)URMN��Sv�&? ���0U�)7������Dr�\���:��L/>X���|;�qr!b�s��f�I�s��%"�h��jэ��`w�;��"�X<4}�|7fV?�_B��my��%1���p&�u�7�'8���TU�u��2��$��5;p�ɝ���M��ES���|g����5�Y��ƙ3�Tq;� ʙ�^Yk]��?�}'���>Y(�ɔ�s{.��O'�}�y)��
�5������*;�_۩,�%I�|��
xcIO�A󪱨����Ӗ7I	 Y���6H7�:"������I6c�_G�8a���e������w��k(�?��W�ՄRb����m%Z����0����uՎ�v���#�h���Re��h�2IP�7s|[�����>Q���X�;HiA��-0]W��		^TIY,A�j��{�JM��{P�t1j�!�rM���Jj<��\�ȶ:˷y�+!hE�M�3���1٧
�jHs3��b�Q�	��Nvv���I�[S��>�G�8{tհ���vK���@��K/ZOZ��0�iG��jP2���	��Y�〡Y�S��)�t,]��U.hAI��^�@�/�%�m8�F����D�+�G�Q4L��m*�y����r��f��
���|�����sF1W�_�T,�[f�ܵ"� R���}S�����\��Bݔw��!Y�������I:�$�����c%8��0�e�qQ�	��$�]N3�
�����娖ۜE��޸k�ee��aO����:	�����<h����|YL�|vT�xa�c�(|ޑԚ����5Qr�ݴ�؏�W�bE6=Vy�_M��$χ�ei���(#�ِ?vØ�͍x��\���C(?2u.o"�v*b E�a�ؘ�.S|�b��~5�5i&a��i���oF@�	=�T-������Ct��~$�u1�����Fֳ��#��8���mD2o-��G�a�͏���,y_�:N�5�5�����x�����ӄ ��׈�Rщ܂F����|��Nu�z����o؈Dh]K�}
�6�ULнL�@g�2��"����~�R��
�v����{2��
aK���~d��L�`���%�۽��`�m��3.���sɂr��*�fxz��J"+�8P�-b�����O�oO^4����I�i�B�m!n�p����0����i0�Ql+���~9����_7�l�6�ݓ+�	Z�0�'T4.�Ɠd�2���lڑ�7Ɛ�w_ϖN�$��o�b?>����@Nt��]c���,���� �X�e����-���B�gwm��\�;(b�Dt��w�}�W��(��XT�D�ař}by~�B.�t:���$Ӭ�U$����[%�������gg�vɮ);^�lGE�7��g�H~��"b�s�֙t/�0M�v��������|�<�P}!lm"⪖�щ�3�AKz#�x��&��NO^���<|�s$��������T��W���1è9�DpU���4�d)E;UY�<9����B�Vz�8����l��?R���%�Tǟ2#F�fa��������FQ<G�����g��*������y���.����Љv�[�~�csk���ud+:3\�#��_�����ꌏ�~qi��s-�'LK�&�]���ҷ��Im��@�����b��c,D�馱�!,X��~h�sJ��׾������n+.X!xK�{�=���;��
�,��ivB�U�mӬ+�����=�t�wD9�L?�Y�~���sc�W�FJ�i�S)O`��&JUG>���_+�D�HK�'�w�Oߴ拔�o��i���`T�K��̔f�uW��=ҁ��0�\B郎d,]Թk��X�QB9����y%�r��R4&&p����q��
�Qy�s	W��p�)��5Q9�n���z#�di\�;~�e���39��@�1�K��Rc��I1>��d��e@�f��:�b��9�o�E���_�\ܾ�t�a�m�^OOK8��{h�T�|� ����m}���90����������i|�Ҷ7��1�c�=�vm�`�����z1uԂ����x����x��5M8�CJ��sG�:g�1Zi%�����V�/1K�[IՒ�mu&Yd�����RZ�XK��mG����K�����tȇ<�|(�aO���A�O��E�#����xQ��e����|>n�����t�gd�v?mYp�����ٱ��)3���w�{�# c��'{qT�w4p����D~��SR3���f�״����E���W ��5�8B��R�.�<�F��x�#a�R"�	�w��
��-A����=��	&��ft�U�`A22��5���s_n*����6}��Y���]���o�#�f�����;�8U>��5�b�z��j��C����*�܈#��W���<;)��u��v��c��s�_U�lf�ƚ��xDG*��,�r���U���{�Ӡ��n��z�7(�GGn�z����p�����}5`��Y�ր��@EЙ/���*�M�,F���n�$w������ǐ���5���5���Q�mC�r�]DK�F}7�yjoqS(a�`_�o}�(�j�`�މ�@T8eCI�[Ey�ڂ�A��쿅2×�L|�+���E�}��p�uŚE�pa�js&R�/9����&c-h.��qA�f~a0�9���\��.�NN�X!H���j�F� 7��z"��q��n��T�0Nf�o��fJ�V�;?~�����
dH�td ��3���D�����U�eӷo�U�e[=�������׹�o[�"��4�0�'�W��Y���'�Ό�G�A�,��J��j儗N �#�Z��Rv�C���"���&]V���	FD!h8����)I.���E;.o(&K�����¶^q���Q;���vv��ڼ�e���r/�P�J�&!��fY���V�`"4���֒#~+ؠ&�s�i*��i���|m��� �I6$�}kh L�ʻI��YJ�]E�~�h�$�{�a���
��粋��U�S�S��ޓ�#Ll��}~V��U���4#f�����)N����w�<wh�.�����k��O
lS1�_.�T
C(.����a��;�*˰��/.���?7��}�L+(&fb��_��r&������`�Űn��N����2��"���S�>]?aml����DV��UA�fT��w3�tM-񸡬������G�3�����,�����"��u
ㅭ�0S1�F���B���ȅ��e�m\8%�+B\vx�M"uF?��ڪ�TM�{�}�L�q~skF�q��f��;�^̝�곛u��.oP`G�`w�	ŷ�<�Q�~�E7ZM[ⴄ���>-����c�O=}KKqm���|O�; 4���Bח���81SMI8餩c��	� {R�Z̲�w��������S*��T�R��"�!㚇w����㜏��K�ɝvQ����>������\t�����S�6UJO��o}�I<Qf�9��K�ܽ6���;�+��3t��{̈́Ҕm��./���{q�Λ�l_g�m�:���$�iu_����C2ȝ}�;i��~�����5��	ė:�dK\MZ[�)�c��q��+���SǨ������֖�|��B!pi'7���^��/��k��;�
��~(`�� e[``�4Y���:Aֈ���X�D�v	x�) �ޢ�sH�R1����q��;��]�?iM�d��F�aP
S�Tz--�n8{�$'r�g���țd�I�W�X�����e���᲎2��� �_"�@	Ŏdmk�ί �	80@u_DK�<z��@�>Y��T�L�}�
��^��������n����r�y���Q���*�� ��1�5uks^N@���ùs=�g$�4=��nh��ѩ�Dc�Ӭ�Y1�_�ڒ㉻��+BѴ�e��
E	����2��^�~{��D���;�	�rZ,tT�����D�L-d�����:�.'�=����O�9Aox��~��觋w�K�i����ҳ�%�]�'��5��ǂ T�����ȵ�ǈ�4*�����>g[�sFZ폻#����m��H�)����-aw�~I�5�܍1��Ğ��C�d���/d��Wr �o� }<�ө��UG;D�����7�q�`���׎�J�Q�@� e0Q���V&��tW٠��Yx9DK���JrGЪp$l��2e
�u��34�$��(��Z�rW�x�V֩s9OW�d���%���xT�jհz6�%gX�W�Uʑ|�J���a���v��%� >s΅���2��^�Vڝ4�(��O�6����͂3��ǼfC��oU^���ǘE��p�XC�B�zqq����'��E0���YK�w�:Ƕ.̝���\P=j��'���=
^��1��0���E��Z:�{�)z;�뫦��<D���U����JN�x�%��e,�8Y-�!�4�{�"��L�#�qd_��L�jp׈j�����r�s�8���p� �d��H��>�i(��b�׊	���`���J��m4N���{2�c��ۢ��
.P�hNj� ��ݭ�4��c��V�_ٲ	��
�i��o�7�]�&˱��!�����>G��Q�-&����L17��a�j���2d�m�b�SU&&X��g��o��r��|;T��FXG�(O�ei��l]������!5��F�
� }h���0�/㈙Af+�(f����-I)Z	�l���%��X�������jK�����|�e��Q>cE��3�� MNX�����@�|6�=.������ >���w��ǡs�'��N�@$�����t4Ӽ�e0K3kw���(v��C�9�wk���s���OK�yE��~3�jF'�u"����q��"����b�W6�'-�ZPN��v��aǝ�>~�P)b�2U��/���� ��%��(����4�H�QZ�d��G?2��M@�ڮ���e4DO��J�������W�!�w֗�ķz�Eu�X&��K�H�}�H;�u<��'��ȓ�
3�����?F0���!�I�x�o\h�=����z׫�LX��^ܚ6�#�7���5D��tE4wR,��ƾ'�����w]�\�������� ݞ-�l�"e�@C�(���D	�%=
;)�{���얂%��焓�3y>�o�ء���"�vZ�R/}}����{�ʁ,=>�;I�N���qd#���2ۮ�K�L��������KϮ�h�Y�Q�to���4�s�0������7(/Z�!t�p���.��@[�@ARj<�t�HGAg9���`q5[���lq3k��|���M��!䊲|/����H�[��6*?{��Z)9N/h	�����e!΀>d��.�!�������n߸7:�r�o]����iSF��u�p*O5Iz��C� M�0 M�>���zjt|`:(ԇ	�;�^Y$�?��cu_5�~&�}S��e!#4��4�¾Z88�mI�=[�`K=j{|����(Y\S�xm<,p���K�B-P	��>!�XD�:���լ�pA�ß>$���k��}Â1r�Myy;�}U�`��h��?������n����W��y��*c�EHy%��I�\�$$��XJ�� ��F����ҳi�d}��.Ct���mz���+=*�|�p�ʗk�6s�d��i�����Y��8p�"ĵ�SD�=�EC|Sɩ��~9�@XNV�k���1P�QiU�'c1=�?#|p��5�	���K��v�>�p��x<Q�U{�{���\��tD�!�riϕ���^�=U^o���SA�x�a5�i�1֧�F���>�� ��f#,�J���r:CS��\*����XL;�uQ�|��:� �Tۨ�2�&��-h��
wǪ=��sDt�܀邳�e9���0B��pV���*�Lמ��¨���KRF[�j��O�KG�}�8��=�����vpa3v�^ZF�PQ�`7�$��n�د@�Ã���1̤!���R@��t�߲j�1�LO=����W5G�{ɖW�^��]&���p��M���X`'�1�\񍡁�A��s��w��4ޣw����e@VA�e/e!�
9�槮��,!T�m�O&p���LW �wJ
�O����x�gǈ�.��N��)3�V�M]��uݾ ����$�����D�"�e
v�`~30Iw|� %`(��FC�~�J�Q��r�Z�m�O)�W_�o�:l�m-��mn:4�Z #�bVUq浭���eS��ϵ��։n LR@$ш���$§��*P�����Nѫ��T����҇���v4+n)�g/E�D����p��w�ļ���k*'�r�Q��LD�������w��j��nb�"5C�W�~�t�_��)��83K�42�Em�,z�QK'ʑ���ƹ�x�x��*�"e|��p�o-V{����9S��[G!a`��KX�����NgI~����,���a��.�y(��xO�YN�K{k��9qE4���L�.�5�)~^?RVSq)Ry:�4�\P��o���H`���p��q��bBˌ�y���V�=�@r�_n�=���=��2�˃<Τ����l�E��k�'ߦ�zfg��k�}!�ߥ���ٽF����k�{��ul�w�N(c���J([����3pj�%n��Oz�c:���D���Ȱ�6F�[��S���Zp-���?��gh���.����^�~�
+[�p�E�1&3VHJ����y�`b�����b
�*[j�W/����ǥZ�1A����o��^̞Q�ز�Cf�}<b�Y������9��w�����%x����{Lʗ�3�R�8�E
��ۣ,Y*! �>z� �0Ro���n���UO���+ݑ�6���5�0˼7@/���S�K|�ۉn�3x֣��ʨ������c*v� 
�Jġ��A�-���.�8�r��1B�i
�����ӨY~��a��@<ĸ#΋�O�Bv~�/-)�~�w捰"�'��f�lt���y�*�Q����"&t���kR'KՃ���Xg��	�����nӹ3OCY�]��F���������!wl��0I��p]"q׫���B}���x|��D�V����-�00J�����x�`��֚F�P��`ߗ� -BN�f�����jL�ē�p^R#P�]b$Eu�G�s}wx��Y#e4�%� 1RuL�����[��ش���vv(E���� �)A���sgKf%N���2O���8RW+�7tS�7�	b�?bE|PQN��MC�m/�1 '6����*�����7�G$��䏷.��l�ĲhJ韐��Y��~�p�D���c~v�՞�^?�yЍ��M{�������~��y>�O�e��q7���؜y�9�"�|z������$MJk�Z��O���U�P5��X���5�=�K�-j!��p�=2�u�zlR!5k X��&.��a8~��ϋo�˫ï��ʉv���IE��=#J}��9,�ߢYRu��,�J�c &=Ek�u����.>��?] љ���bP��S��Ě��f������+uz�޳��(0�z_�";�0S�����+l���D[�ٿU������U/��2���nm��P;��_bK��!��Y_i�q�V4� � �Y�}�0��Qq��<��. �wKK����@ [��::����`�o�үKyH����q�>�)j̳��Π��q��p����x8�l>�P��a���?Ǉ_=X\e���#�m*�X�\	�7�~Q����dS��a��.�ME�mʛ�S�,>����|y�!,J���+��w�r�!yCu�Nɇu�qp�	�!J[-&�7�4pDR�~eH�g��h�E7p#��z�j +�!1��f�uI������	P�&�-zߒiW��g��_'�	?���_�����!�z´`͍i$)Vl�JeP�q]yt���`�݂[G<�q�q}]�jK*.,NP��6���s1�{�Qj6���:7H��nQ|��J�[���QpC��#�L&�v/�f�g��1:�i�zn�Lr����Ň ���%μo��v2��Y�*����oǘѤ)�� )N7w�7�h+�IP.2�zzw� �L�G�|9��L��ͷ~��[%y~ ��S��Q��ʿ��є-EFy�y�?����{̫�?q�v�w��J��8��$�9�l����2��M�<_U��\K%��s�i�1f�� �M�g�+R�����U HÄq蓥p�y�f��Co�6C�G��UR����V���(�~>H*���$�˛���j����M]�M���a���h�4ʀJ�@������uZ����	�� Q�'�4o�S�s-h����/1 �8�UǏ�;�k\����b	ŉ:���`ɪ���Q>4���`7�僗��Ҏ��$L���ڵ���@|�~r,����>�.|ʏef)�m)��h�
���*�Ԗç�]6��D�I��Ҩd��242ؾܨ������̘��Mt�a>y��w���A/66�$�dN�&�����b��6�{:b	G�~�ܦQ�m����|%���0d�O������Ѧ����M-�C�/��.K7l����83[6���d�)վ��A�m�A��Ō����m�*OO��D ������ۆ�|{�(��j���VCԠ#��B�B8�"7;��1����XC�J����g�(4ٮ"5���|ib��K�=H�b�A5�'���J�F�+���1fm�w��Y�l[i�}���a�Od���D�ȀR��v���똰��u73d�9�n��7� ���]��D�t�<f�3�mѾ����(��8H���� $��+wB�1d��9y���]bK��Q҂�U{L9VTwxhyӺ�ct�R˻��ر���p� xV�]��S��h-�S��7���n�6�� 4C��O+� =��I��"��$�4�[;V�mr��'#�-M�P�w��5� rz��јz�Z\�;yPXz/�a��JPN���T���(�CC�n��傳����! S��@�>k��)������N��
Wo�
ɷxF�N�k����/�����Qc���4�����7]9������[�����,"JÅS�����WRF��=�Ltv��`&�Tl9kvv��B��'0���b���T� ��d����t��X����>*O��r	D�����Ǿ0Y� ލo�rF�-�����=^����X���AU�\@7{�BWXuYX��\r4�w�.��ߗ��M#��bL�ƣ���H.��ѫ�^����c�0(H��;� 4���Ĉ�A��~m)n�8�kᔭyq�|��J�`���7C�<g��)o�!���_�F(���7��Q���[F_�f��@�c��1�1jqK�R���kM8�:���>cO�n⡀%�0U��'��ڀb����̝9
��_�L�g��R ��$�v9��U��Q{���+{�WM�6$k���#���n"YH2 �5}Ĵ��IU��5�H�p�ݺĢEHGrs����}���4��!�P����-�����6�r	O4���S�-��)�jက��oa�V,�[9���/R|���2�'/g��,u��r�b����쮛ߠ�����qk�b�8�}|��}��_<d�
m���)K�F�0	!�d6@��
`�qC�B��n{�%d[�����͝���G��0�
X���y�Qħ���rlw�=%�M�u�՚�I\k^���y=�0�2�(�-�- 0�� ��IC�o�������x�c�L����;�x%�?�״�b�@��Z �
VY����2�'c����UMs˖����hW�uK��[�;���G����$lh�l�Z��ޢ6!�@ŒY��Ƿ�C��i�#SN�x���_y,h3��jc��Q+@ҡG�pA�$�m��� ���*}[�5�|Uʽ����z��K�9�m6�I���p�j���?B�+�vpw2:�CU�� Z��@�� ��[��Ԇ�}��"�f�`}b���c��#7�1��'���_d4���%�`����3��� �R%%L�U��E��Y2�W��Fh#Z��R�1RP�m�8W���¯�|�=��G��xT�H����q���J�L!��U�x�Ɖѥ�\��sm�2$�'�"� ��qms���|�P*u�Y&o�P��e�:EG$�iZ��ո%Gj�Bn�Ⱦ Jb�)wDr%|G��|E>�vDO�3��0�{Fs��[���eu�Y�#ZBLAcG�A�ydlZfe3>H�s<sث�I��p�.�������_���boP[�bbq�!�겪��êB:(��CF�B+\\VFU&��:���9�[�.L4���J\�C�g0M�����1%�*-S^N�u�$��^�}��a3�Լ(�6n�b�3�-��lf��j9�񄤲�I��
�}���Q�vM"� �w2`����n@%\b�M����0�<^ڽ���!�B`sσm�M��Zj�����ߗ9�"	�����SL��ʲ˰�`b����6��Új+��(�ꪴ	l�H��p�gK�-N�,c�mA��em��B���.�IA�M?�>k�	e7�P+�[*\W�ƻ�5�����$�&H�wN�Pb.�x[:"؋N�@?����m���ؼHMHy�*��9��6y*$=��)k ��0S��1(t}�z���\�7j'�+1��r�~#�x��L+�̎)�C���f���Kz�v.z�!F�:� ̸�<��L����]`\�'z��u_��D�0[�E�G��J k����V:?�O�����OfoʊG"�b�HQ'�Ё�BK�H�u�jֹ�V�C�n��*��P�EÔjB-��z�Ё�|Lc��8:E�I�~J1���::(z���~{�rtSx����&z�*L����E���r0�J�O)|2�V2'qʀ}�O#�xF*�x�|綽5�cK���+��'{8>��9��i�^�i��iN����tA��!���S�-�z�(���V`u\`��7-�F$E0JC��cbQ:��@��n���܃����k�P�#b�8%r�\A��<��oொ-ȥ��^ͳ柀����ڧk�P[������y����M��Q5�t�Q�j\���3y��oq�D��g](�G4*�&�J<Vn��Y��a=D�g2+��H^腏��]��gF<�Ji �b��n�$��^�,�rP8?4�h����(�-�L�[B�T�@ZE�4���M��3����F�O|�Tc���Sw�U�����e�8MlPȷg'�0ko}�ŰͻDz�.�zR����as���=�]U�6%A�&ek	,�w�\;�m�*<���Q|��>G2��}VnQ�W��.�u���v��3+�C-ݼ�g�3�2J6N]S��B��j��ǴR�U���._(�_ۡxǪ�<�qt�:�B≟�=Z��a��ݻ^�  ��Ӳ��+��<5������V��r�g>
�T�/��ϷlgI��z0抮:�~]��z�_���8A!%�8WNkd���b��j�6�{�+{�[%;@�z�'`����-��7���e�e��	[�����YU(�%�M Č6K��s�R;Ó�2s���V�{�vj�'7)��/���Ea�]�s�/V(l��G�~�i�����<N��,���c�n�a�.1��H��;F�r�j��;fH�[�]�^�="��7IhI�RؗG�7]�Fl��8�νpo� ��7�.�mɉ��0ݤ����Ì��0�2[��{�?!
�0����	u`��4�ϧ��������Q�#MJR���.;/���˶9Up�#�^��D��j�89,�O��nf� ���������g�_�mz��3�o'p�&D�Tz%�Je�~ �����+zF��fއ��J�֖���Tlr�J&U�7¦��zDg�#I����p���*�?E�U�_��J�Q$R��c��X:�cO�0c1�x��U����6|���üy~��=���#�v:Uޓ�ה�TO_�H�SX	A�^���L�o��R��'�3ﶍ)7�D�Zg~�L9����o���2a"ہ��x���H<���=���]ᗖT?�KX��s��2���M��T1�dUo���D�!�E���4���ZJ�LYg��y�V�E������'�!Ҕ��[b'��z_�%BT[8>�����T�B}w-����ؕ<7l(�/�;|��D�l�z�q"	.�A*6rh��\�&�@-�P�,�>NX�^�"��)տӲ>�<�r<���)�j���xX���#u���7��^��m[K�daߐ�6��Q�&���Z��i"�l�^�1$��%��I[)}|��;�8�k+��!��R
-��E�,��/�07M.=<�#���i�f�R�6���2O��M��j�A����D~	i��&d��U�� �W޿�pm���_�+=p�Z�&�(H=2}!��q����%�����{T#��W��*j�H,�Z��m�B��k�t9)Z����SV�u&0�rh�G�ܲuh�ȼ��n�j���ķp��;�ݍh��sJ�G�\p�]J9*㫵���g�6Q�,A{P��=~L���"�{���n]4'In�w��s�ǻ��]2�X<��_\�ݫ���e{ޣ���6����<��r&��JUL��q ��fu�b��ßL0�1��dM�w'��%�H�t��󪻥�d����9rH���^���z0����&ڪ�l��%�Ƹ��U��Z$��T�R��k��<[_����^"�{�j�X)4���A�`s胜��6��O��6���\v�;S�\�%"��0���$��%/������jN�-�訴UY4�
�t|ӂ���_�	�Ƥ7>k��c��F�Ǿ����*;�����y�U~�ǜG�N|�š4�V�n$��.�N�/��CojUj-9��� ����v�ၿ����{�Q.���	<|�u������X9�������#�&���z��i�A,�  =��tq3EE_��F��9�+�N�iY�Ѣ���G=��م��ۓ5,�t�"�]��.��LU��p��"�x\@Af�dyL̔�o\��v�蔍7��F���gD��-�|�>�Q�>�p�����Y��I�+a��/��(cR� �}��l��R�<I�f�N�[d6���nc��Ghj�$9�r��!zc�ɶZ]GI��eN�{�p�<�Qyz�?���eL[t�*9��4�?�c�5�D15�$s��cU�Mר"�dD��w����U�U}%@EB/MFA�w ��DAI=�+i��kg�����5��R6���n�D���ma Јޚ��A�_�#���9S����ȵ�m�ʹ,�+Cr�N�ѪA"�\����=�>��ܑ�{��&=�k�?�����+h��\a7?��/Xg�]�����{��\؇:t	,ª��#������~�$��������[e��&ļ L��#�J�{?z���U�2MK��5�p�;Hs��'`��jf6z�j��9(�l��F]���NY���ҫ<ه��_��k>�=�V��"���Ỳ �[�����Zi[���n����!���E�Dx�42����b�T���������<�?YX=�X|�E�u=?���R�s	߮��.�Da�(����W�S�f�)�~�w���5�� �߉ `��݁�EĞ�,�b��#�?��e�g��w�N��-|�K�3?������(�z�*a$�y4|3JF�>B�\vN[�V��'#��m���S���]<{j/��7:N���:)�m�I�+l'���ǩ�\t8�)]�����p��lX9��o�u��J /���,��� k�&h�P�j��g��<H��9^d�6<ko�h�j�>6֡�e���d+�'d���7%L9`��p�+RȎ�sXKI�A=���q�܂x���t�����Z���H8'B9W����P��uj���$C�в�q�{���k�G�o&��K�2����裤����O)�X��_֛U��P^O����|�M��\�L��O��	�2Ml���*�)�П/0#�RjϚa >nY�~ט.��[���H�"VĀ��\N�r�� � \见̜��u[�85��S.����S*`B���8I�t��pw#��ឳo���}	�>�8R�Cv8n�D3�Z�b�*�1y�LDx���y�:�2Dھ����)��������Dc���&&������1�&,Y$�ah3�f����yҞ�q��?�"���c.Z��c�i�U��NZӹ�I��)��q\bӶ��}�����\X��.a�b"�\k��*n� �+�C���M��$��e	&�C@�P� �����)��
��*:��F����X���}�rE�S$���"ϩ�
_�`N_")6��nݯ]��Q�7�z�����N�,r�z��A�� �v+�^������vw��=)�X��j�R��̧��3˙¶�˕b��Y�я���4���2�����upN�g47���猡��oc4sG��h�N(Lա�>e�/3����:����>.Kz{����\��﵁����Ք0K�r�0Gp�%L��w�2��{X7Q����x��y���GHe\P�s�p��~�l/q{����4A�>�Gm3�G=��O*�����e���.�����a�v+He�����o���}� ��uV�GC�@b$�}�U��@:��["ᐝ��$)ɠަj\+6��	��pC��p*䲁�x��F�j��Nt��s�^c�p��U�%��#�I���<��P�EB�H�O:'�<:��@HSfI/�.��Җ	%$��:�1�Ԣ�`{>>�֫辑�dI���o�b���	{�=&,�D��DF�]�C��`�*rŲH�[G�}.�h�k^����_1��S	?C[�I��n�	Qh���D%�Vp�M��I��Q51:x#���ٚ- �m=�&Ξl�K�k��;0U�+V�>���]C�b��Ƕ>f+��cu�ICؽ[����Y$����!z����!`�Z?�?D�8|��r}iQ����)%�9��P�����(��j��J�+�'g�$�lJs���*��
� ���1s{>����o��(�r��V�#5��IS��K�bF	��X��V�
kW�i��8�?�;����$N�4(��^�Vh֋!mҕd24	�h�C��V��I�?fwf،�VO]j�'f���_�����d��R�${��\4
��'�:�o���xQ�\#���g�Հ�i����G��A��lE��E|a�L��W��&j.w���(z�خ��0�rf�s0�@_�."�	(�Ԯr���������B�'�Iu��V�]��֌�F 'O]o�#�HYv�Ј�7��`垓`Y��_s������1�W�R)x]R���͡�Y$3$��:<�X\�<�������/Xr�q\�b5�7]�zEG!V��Z�v3x�5�rR��2�~�6l^�O��w���Z�83��FB>h��HI�.�����Z��P��>����>~�zP�:�{�i�B�1W�"��_��*a���"0���`p'�9�k~^��h��h�%�C�lQ�ܫ9���	��v4�&:'d���CE���M+�fkn��H���6^v��-�T~�ܘ�g�';�*f��i�#f�����6�K�]�2;������%��#� ~Y�� ���r����A)v6�����y�pG4�6j?��fM��yw�	��m}�.��⾘|\���uy�JEҰ���*������Fy�e3�@:��2g����k�{&�a�����H��G��������ו9��A�`�Z���]�25����/�7�V������cHl٫6jzo����8���h�WJ��W6d��>z��%�^wm���!鏅�����f�*!��Z �#mE�l�<�;")���Fz=�������\YU���|E0�9LlƩ/�{<XSOekg�A�m�f���,�����o��m��ߣ���,o���oE�I@y]	k���t
}���\�KKk��1�V�=Ƒ%W`}�ow��3�
��_�kp�A���	�����W2�F�B�y������zPr/�=Wd���~���mH�2$��O���+y���t4���`�a�EiO��iܟ��C{�Q�g[i�:��h�I^t��M�-[��K����Lr�D��O��<NW;�Қ��jf�x�IX(�W�G)�`U�F�����܆�hꑫ�����P{6�ٻ�ڗ[�q[(=���+�ѐe�f������8�;��h䬱��_�=�>��O� .@���3�ӵ��	4��d���D��z�m>4�坆ir��b:�[�h��Y��X�Ӣ���,;���BA��@�Y}��=�p��B}ڏ���R�3��0��0ؘw���<՛,w��Bx�{��L�Q��#q�>�H� ���ȉ��0�m���>�4*&������-C�x�X��j�o�X�B� m��~!w_��Ys@u�6|0�2*(��
}"�֟@H�.c[�¢������ �����h��r^'��~��F��d��Ĭ��"$�.D�Z���l��Ql�I����?!����tI{9��߉��b���K�=�n��`f�f�{�,�%&��5b��U��1 |��� (Eڹ�Ǉ��c(x">r��N�C��2Ӷn.F�5��(��}�����C}c�V���GF�x��Z��TÄ�ڱ��춘p���s���čbg�!�=2V��M,��$^���`u�yzz��`b��/K_rXGj��9�GV,��U���Ct�Z���rcey,; �O�*$���LѮ*�\���#@����.���	�iػL�ѥ3��Q�q]�1=��-�07�X��2��T�u�ZQ�`�Ɏ�i�\��@Ҩըs�0!6����N��i���}!�bA<�Nܿ@���<*Ӌ,6cQ�=~�Un�ߕ�'�z�Q7l�7��`H��� L]J�%jc�?3��ko��[���7h��L�a����+�㽈�l|���ڿ�_Q��@_�tc���ht��\�i�_�xF,���j�O5��4hJ�L �R;/يp��NO
(�j���WL ����۠�-�$��;n�2;��kF�uh�qC��̝4n�5�QY�,�^���F��{�J& 6A�M0-�[�c���dG���������b����FV�nw�7"Yr.���03�޷pT��ۯ� �2�I'p5�n����'T0I�U��=J:���6)o����衟Ac0*Q����F#dL!��F�7�c�!u;�2R��T:Hl�
Ե�'���h�)�:�i�s3�|){���9��D�K���V����dx��\�������_�L�.<+���{�������{�[EE���tNR��J���<��a͞>�J1P		Ue� � �`BA��l}�a{�cP�����ĺU�����d,��[� �%.j�W���*�4���Dp�����^�T��6�H�)�oN�<!p��D�m�q����V��{$�{
7�\�|˸�? lw4}E��z��)pH��R8^��ژ��8V-|��>4�iξSW�f�X��60�$�V����h��v�^/�><��`�gP��yu��qa\�!Cv�H$r�Ӑ<qe|�x�±w޸�X���X�b�M�G9��y�hI�T]���0��~{�F4ee΍Z��W
=9�b�>��}��p��Q��St���d������4A�Ѐ���:�c��+~]�R�A����x�-X�T>-5���_��]!�SdF8J\������"9�0:r���EA�F��Cb�Z����v[Sz�[+��#,	�A�^�<�Q�E�ٳ�6�,�UU��O�T,����xC���$��q�B���OA^�Ԅ����t,bB!P���[����a�T>Ә���l"U;�sK�TO����k)#���

;/�{� <gq�-j�B!.�tj�%�ɯ�}Rf���Kuݬݣo��(��aC�@�Y�c��>�3#���	�jH���D�Bє��'�Z�j�iN���t%���0zi*�;F��s?�W��={XU���F�,
�G��ո���M4(<���a�a�y��ZM����o}3��?��-�9��C�z�!H�A�YH=w�Z�$�c �be�ؐ�A��m���f� {N��L��Gd�D�Qe�!��[���}��Ǒ�X�6��wa�
�3�-�%�9]1�x�3���(��T㈀���Y؈�vp�m�:�y� �t�N�>�,,c�i}��]����c�f=*�	b֦����i�^����1w�K� �i#0I��La��zS6q�1��0ĺ�C:뇖��'�[56�N�|��3%����^?Mp�-�'IG���/�{�,����/�U;q�*b����n9���0aP_� @a���#�\�q�x�kKGM�\\�gV�~Sj�������$��"�@������H�(#�)�&�x��`N�٫ɹ��}�	��C�f�_���/��r����F�O��1�|ȗs����ы��R~0KC�_ex�x��k�i&V�S|H-��v��g��� �aNN0��tQU�{�^ܶ���\8?v_�Bv��!��]���E�w�F�z20�@ǩ{�0B{D�,�=/�; 7�K�b�������YB&�rc�7�}w�NC�ߛ|ը[�H��7� sۢK�g�ӃU�@�=��ӻ��h�g����4���LwD�"�E]�g�;��TE�E7�EC�HdA������:�X.mx��|#��	�#��mi+Vn���y�8�"txQ�h@Tc>�Tȧ�������v�(���FU���Z>pC-/h��!�����`\~l��w�>s~�]K��ru�$�V�gyuo�����)���<�@���Naĕ{V6��F������RGo.f|P��1�N�	�A S���іl�?��h��P�Dk��	����tv7�q����D4*h/<�y����qN!⏲o�a�7���%��!p��=O�䑡Y�&F0u���Q; �Q��'3l��ⶦ$JN"|HT�pQ;*��R������wd��Y�_r����}���A��zQu�F�x ����}��N��$���*9�Ij�j�	Er��Zo;!�ɠ��R�b�B?R��t��99[���`�;�g�|��/@Sw�Ȼ���j[+�!���}��}���J�	��a,>������p�{�(ɥ�⦤���H��NX>ן�J �uѫ?�N���P_#��:%��P��)g��CkB��\7�VT}K���:}T���|�!��v�$����4���K;��I��� p�&򢜓H|jq_y�O� 6�I;��[>ύ$��m@�&5��(�-1��ڀ����	av m+�>���)�a�+�k8r����X����C]j�ی��<�W����,S������Τ��׹p�bQ��s�C�+V�-D$�*AGݻ/#�o��&��Q(�#�>����L��E�d�����y�����o����Ȧ���h�Y�١޲j�歟�O
iO��k�<$}��Z:W����[��9��îF��]�*�T�@5B2j�R��&������(��%�YVo*�7���~�3;t5Gk��7��­��k}�1�B94�o8Ƥ���л+��l/e�R�h�m�Kf�V�*<��g@/� ]�8%b��D��j�d]�_�;���ޞ|t�'�,�>rp��1�0˓��Bi��hF�rx�$�ePǍ,� \�Ve;��J��~��$-	�b�"��H�+�kя��-�G�/5C�rvxZW)T�1�� ]���
�>���#G��*Vx�I-c	�#�n� q��*�T�~'#��%�Ǚž��\<`��K�&��ߖ6��D�)&NR )�KǷ������z"���Q�mS	���t\��.����{�]S�#�*p�!x%| )��SMpl�E9MV���nq�W�I��a��,?X�f�5���5��E�b #c�a�������n���z��`�0����ӾD)�B���;@�;���key�(��f�m!��9�6���-�i\����Xǉ�[��e/��t, �U��$�g���Oa��!n�|P��ЋX޻xc{Ȋj�����'gy%8k�:���muNU#�t�}J�ܙ��`�6��!�m��˩aq'2ɨ��W�1����y���'Ӛ�H�3U0�#5�푪g!=_Itiw�UV?�b�W�d�Lz�G*�Ef���M�#K�ޢ��N���0-��ɫd{/,����y�x���RO�&��G\^o[��+�_�In�R���*�Z�[w3�	��]�k(�����~SG䭓��2�2�[>���g4�\�
�E,��/�);B�͝���VI���B	��D �5�+��n���LG�m�?8q��ܷ���a�~{c"P�Sw{#m�h�7#���$�̺��L�j4�à�e�q�U�]Z�.cZ�866#R�пN�`�"�{Oh&���1��D%n�9!���e�h� �l85��Q�iT9Ȁ���;��>���l�53�����IQ0_��Ry��\�ӄK'D�K��S"��	�ϳ��t��L�f}>����c�@�4��vO�i)P�a���&����3���b�T��O5���6�=��L�R+>b�Uj�e;F`6{���AaG���Rm�3�� �[�������ڍ���^�x�ne���1��Zu����dv����D����G6��t�Ȁ�+UW���Ryyg����K)q�VuǛ��o�F������0��M�>��������n�K�еk���SC[�t���=�m +�I���`ͅyTBM����	;h��h=��<����DR�"����7�^�Y�spP�<ac3���U���w�e{���Z�
���	M�w5F�ppfJaW�~���ү��D�C7s���?F	و��h������
��\6��Hw����'��1P�N}�ӴN��P�Ζ�"�[g�<�H^�ć'�,���V}���k}������~�+ª"9�v�=��$I�N��P.ީ�e�e#!�(/������L��*��Y*��[Q�zO��c�g����`�{�&-����A5efA�ek���V���N*kٖk���"�Gvk?�����{��W��J�D��?Q>ٔ�=��ᒒ
��Uh']��������c]�;�獪1�AI@E��&3�a;C�Aq�{ 6@4#s���W>&<q��xh
u��(���jl�ޢV۲�c��E�t�|�>��R�߆p�o����?��y�ܬdr�c�*l��B�L�"���t�!�XD�\N�Ro����q}�qx'�/�y�Zfx�-4tC7����o�8�Q"�a�;�L[��'
(�Өmj��0�*l��D�aR�ew$9i�0���A�0�_͔�P��U���\E�\i-F3F%�}ˈ��7�~$$�E�Q���ޞ�.�=$��s��g���*��Qr�����Zη=��<�pG�\���Ų�3J?A�м�ES�mA��4!~�Fy�kǻ@�6��u�	��NT��n�&y\|ER_=-��m�,,_�#B_��v u=)�ָ�����F3l�>%����2É��ؓ2yw.*��ꍩ ��V�nc����'�������
�R)AG�C�&�ȑ��ǌa3��G�u��1�wT�3��������6P$wa�6ƛ�"cc������LPx#��h��m�������V�M1�u>8i�U�N��Cg��S8���Ƹ��@DC���_*���4t��#��U�T���DGTj��a#?T{�Vyᭂ���?�#���M���aj�����5Ú��֜ks ���y���]P,��|�6�>A6!tn]�õ�b���N�T��/5J�ɰ�\g�$����}t�kװ�ck�t�4��d�&	�{&&y-R#��q 鶭��eNB%����k��u�`md=��%K展A�$?�N�G��s��,^��ΥmPf�2!��.l�n=��U�����Ek|p+X��cϝ#�l��/�LD�L'��J����2h�7�E�B�0��Z%39K�R�-��b��o�Z^���*�d�3�(���*��k��0�0�B�G��Zk�W{J�3^��2�H��94��'��ݒ�a��n�;�*��y�eLO���㵢�:����E����Q�V��0���77�޼#�����XJݚ�;'s�S��,hDP��:*��!m��G�]`ƛ^\'L����W�7�:�=�u�[�o����Go �^�P��%0��I���^��^���:�^&Dd6`mp��eb��=��A���;P�C����
�o�U�L�Xu�<_	2�ikL��u���B�Q
_�m 1�~rj�Z���@p\�@4��d�<����?Ck�b��}��`���Md�b�g��G��e��d�ٵ�����8��1�$dT@��ʔ���:�{��[(f�{C Z�43�D��m>�$T�%�L�adw\��6m ���LD@���2�?�}��m��� %��<&_�ʤ�#΍��@�ڔ-���3�|o���̪tAG��lI<�%��#��3�C��;�G�^���?	G�tms���H%=�F��s�!�-D���Z��{���"b��6����(o���:��o�n�-o�����B���6�_Ϛ ��
㻥�s��%����.�<�
	�+�e�"R�.�J���v��E�7}iτ�������QQSu������9�)��
�`M��|]�VV<��#��2��i���^�d-yd�F��p��An�����[�F��C8@i��=�t��d�ڙ����'C��}���q�����l�~���h�gܞSi�Ϸ�&E�w�/�!TV�E&~��G<�hJhʣ���*�)�|���e��+�*�Tl��=����ң8H\�1��{���1r�xBiz�������J�Y\�(xM<bp�yW
��m\.���^�X�Oq; ������ �����Ql��8~o�W��V� �=�YR�X4>�	�۪8��b/��N���?�}����}C;�s��^8I0�c(y�r�d�	��؞5��_��O}FWG�hq䎭�r�[��=Gi/�f�@�鈑�}�Hi�i�#]=�h�B��A�?�6H*�YG�w�RZ0P��5�{۞���uX	�5	�%��`h\$���c�q������x��]��`Gz�0�3�E��a�'b�\[��{�C��
ZR*v_�؈�����y_�03l,�Ky����t{��Y�Q��
!��2e1�4���ŀ"��V����H��@I�-䫹q@lɖ!��t��M�!4��`�R4���Ȅ���=�~?�y��x��*�@�%��L��~07ZȢz�I\I�_nZ��D�k��Q53:d1�a��x��/Y��;��r�{|���S_#����l(gM��N�u��GEľJ�	�����)�u,:�=�o&]��:�NU�k��x*
 &�nƃާ~=��/ڍ��n�Y#�؋po���v7͟n�.�`��D��h̨�}ƃ��4��89�J�Xb�S݉�����'�X|�?�����!Y�N���dЀChb���œ���ɶ������s����<Ȱ�/
��>g 	�Sͥs��iS���55H�Lc�����A�w}Pn��,�[(�Ԥ1]�o�/�P���,�M��~�*�4�㟸XK�<4+K%�L�UTZ���g.�#&�Z�cm�e�a|�|��Յ�A�A{�1�H����/����O�'�]�hL)�������O�XώkN��ԥ9�jh� Nn�@CYL��ߩȸbQA�)���*� t�!51 hYL�>�s-k1����x��htc8:�x���a�����F��<��K zQ��u**�ΥwjYЩ+�!����|�C��|*�����0F�3��/`ԏêKb���lmH�rVP�%�Z9N�:��W�/ȹ���N���[�.�52;�oH3{I�5<�z޸�l=��
4�Ӻ��G�K,.��������&i�)��K�����z��kK$)���\�$6oL��́�l.>T��d�}Ej� ��_4��MкH�t��6r�
z�hF)T�:��/�A�h@���С��f�~m�N�Ǎ��t�^���wgZ�o��}⭁8ϖ���iXc�fP{�[o����Bu\i}2�7i�2i!rP�h;ͫ�(9����[Q�)���[���� ��ˉ��=�Wn]i0��W(���l ���-��+�� _D�;��-�1�S�����j)� ����U��GH����G1=�t��Q1��BSw.�z��L�W��rY.�~�3ڌ������e
������?��!S��~�
g+�L�L^bo��<��H
���_��YՌ��I�T����vG�7Ua�.3wp4���d\�!'6�y�0��?,Zo4�͈=��K��#�r�ߍ�&1N���Xr��,_r���J�>CG�Y�?��C~.%�^��Êc�X�o��= ����-��� #�u�]hqF_K���<�
�W�J��UDzBf���zY�0N�	�zG��b�.	��W��w�[��΀Kx�S�1N\�O<�rD=�兖|�L��. �*��c�׊�Ժ��B��&G�a�޹9����#1O����I�X�%�`Tm\Q�f-4��eC,C���8�ͮc8ʒ�T a`�m�ʇT)�ס\�ΰ�U��Y�ˡjvH��mG�=r�IV���'w4�R��αR�����Rn�r/�	)̢��i�����B����i��E���򯐄�e6���M� ������B��b�D�����唓��(h��x,w�˭��b_i(���5.R.B�И�����-�:-����ֺ�gC��M E��́�u�v!�6�k��W�P�#q��^�z'�<S"�A�DM]ޏ֚U��",��T����<�!�[H�?���_�e��|�%� [m��P �\X����iϣ)��*p"�-���.��^_.���$��������ck.��e�A�BM,]1;�|�;X�DE����h֔4�e�s�A��":�*(V���Ч��/�m� d�v4{��[����p"[,��i�-(��i�hۧЂ���Z7`���Y��&����2��_t�"C�j*��H���DE
cY$�����-�g��a(-���g����(	:b��A/C�W�X�/'��c>h��\�r�՘-C��*)��6a_&�`��a�"�ԯ�5m�o��\.6],P�a���T.]Œ�7F� {ea����ެ�.�/��<���L�z�
-���Q�s���ޙ'J	�]��ퟥX�~)���m�v�m�߇B�>_~ȟ�i����/��\c3�}TR��u�����w�^�\%�����[��$^�)&��	�~$�l�J�pxBd���ѭ�f� ;*X,8�eB���{�����=�ʮ_ȧ���l�Jc�� �|��Y��T�Sg����PC�W}���G{��+u�S��g?;�*�����|h��E�l���Z�����E}�5
�� ����q�H�鐃��.�_��O����C��b�R;y��oݨQ�1;���p��o�E���0�9�@�����Y@3��g�[y�$̿Ț@��zns�lϢeVu�$̓�?�aN�/�B_��e�@�E1K�'�)���gh\�p~��'�@�ʳc ������+�/�^+߈H�Z\�ET�:�r�ӏ�r�/eMz�Km�X���|����`	��^ap}0�Z�Igw�����}��EK��D����$�A�HZl�Fu�w�'�1���"�}q�L�r
�bX�6:I1{cq���������. �?S�����pY�!�3��ڃ�����0��?�"&��CvWz],�I].�HKt�[r"�	���	�W���Y���dI���T���_�z]1Y�?�P���3��>��\t���s�$0uH>�;��&n*�w�Y҃�FBB�h��h�{X�[hK��'oFh3/�n�RL�Qi�jܚ���0ν�72M(W�"����/���:��6q�dr�٩=�#�7d���D#��懕q�a���#�m_a韂&��9�����fF��:���c�����H%?��OpwcĨՀ�ц�A�^7�Wx���C�D�.���qF\>��,X^C1 `ۧ��MF�|�����Q�� C�j�a����:��`wۣO�y��xj��q�NB�	�d�����T������?'+�4�2���V�o@�d�78�v����s.R�����?��4�5���?&�җ�Sx����*�L�1��^�+|kؿ٣�_�ΑۛT��~��t�`����*��p�YT����L�Zܔ9	��#𻸋H�aBh��2�Y��P�:����usI`�*7�@����&��`�,���>��՛�������L�ڸd�"���-~8Z�uw��	*0^�<]s���	JU��#ZHv�)�|Q�IL����$(G� ���A���J���]�:�:�s��@¤Q����ub@a��m�9>�ײ~8��`�͐K�K!9�]G���(��v��"l�K����5s�� ����}"�`�i8��Q:����)�j^��q�����7j�o��{����j�	�C����0`t�D����w��(u�V����;˶E�6�Ͽ�$t�FiF�8Ģ=��Ȁ5���Tq�յ��fˬN"q-�Z���)Z�&��Y�b��s�B=KQ��~DZK�:[�oc뒚t�_��EM2Sc��=l��<�ɫ#뒑e���~u6BA�#�SEg��Pۜ���pǙ�a�q��w��\�ާ삍�U�[C#3�b:�h��K�yG����@����O;zz��
�f~j�͕=a�ES��p�<sΜ__h[����hUZ>/�lk]���H�u���K �FFfq�(�E��)���u$����s���B/3*�8��8�ޠ���Id\jT�0��v^*���d>[V"V��ep�p�)������a�-H�cKQ
�zhot0�B��q7��i��� cΑ�C����fDx.�Υ:$��>����T-͍$}��('cC�;^��Ck������V��]��zϧ�0�v=6��q��b7������I]x�W�_o�����6W�B�%��C��	P�����ձYZ...Q>^R�� ���������a���4�s��xE!��gbGH�Szu�j�2�(��������x�.r엏���U��LO�,ݠ����E��PI�浖?j�@��X%��YN��C�P	~7f�\������O:����3�X���rI�.H���Y�k������#���$�%�*a�^E�(KKQ#K���vqޖ�e��2�N�A�8q�D(�����?G�(���!{t4�hr3�t���t��NV�r��g�3�4�P��v$�G1�h�vD�ص"�٭��H%��5�qB%�*B��To���)!n5>L��L9�0DzL�)��9�@M�}��?L���dە1sz��ȯx�>�a4C!׻���ƒσq�t��M�Fv.i�=����+i1�vr���F�t%�������s?���iɄ�f\(�j������{��F%?XG2>j����|��aM�z���o9t��dR�]#���^q*���7����(�⻖*��̚��6G�WMI��[�/�"����;Y^Λ��ݣu�ٰ��B��/��vZ_�0݃*C��j+Is�`�pӇ���YY-��4,`C=ä�Ij��:��޻���1�\f�"E�6�٫�;V���_�Bh�����W��\+9�����ȓ߭�h�!!��'h��:���R���O����\��n4r{�G�]feE���X�AK���R�cq�Q�'+�	RK'Yǡ��n��7 S�0N�����q��)�8�C#�a��yV�t��t�n��	���O�{�)RK���@�!�q��C����Z�J^q�y��r��h2���f�	�yA��!�]�QL/dkaǆ�"m}Z���0���������K6����TI�[��k��/�6�0Z<�l���2a� �j�ϩ�!=��� �x�Nl�����Q%��.yt�/3�=0�zGH[�Z]d�[@ݮ=�C�]�kfЋ�:��Y�a�0_{	�Aն�����
���px�Z?-�I�dw���XU��s����96�	9�E#�Y�VG�����{i0�vճ���`7����l�A�h'o���4���m���*��0i˨�}�n?���Yp��8�;�m(H_1��>G�r�\��ѷ1�1�Ȟ��Ǉ�"[z�:�2 �2��.
ij��~7���x�LӖ��nnޒ2�u1h@qH�X���fdJ
^3>.�%x}���"���Ҭx��5Nw�-���U��X���ۊ����O�Wp#�:ߑrN���'�4�Q��/X-�C	)��@T�����ɯ�˲��%èP�r$J#LF"y��^	�:�'���U=~�]���u��3��i����Fu�`��ǩ���"�S��Gn{���ċ�聉�ه$�V��B;5���{<���3$�_^���>.`�<��f��S�ԍ0A��t>�e�Ћ8�d������|��7`eYy���o�3��x�(»'Or�.)��M�ƽ7혳~��`���QKc�Ŗ;�z;g����<��k�o�gφ�2�*�r>��s�do�ϻoq=o6ӝV�7'l$@`hRc��Cƅq8��*m������RIjEUw_��M#��B��-4��4v��հ�d�xJ�ɔ�{������������Wظ�����J?ϡ�s��q��M��08Ow�w�'�0�٧�~z�n��_N
�n��C�����Q�b�Ń�ml�D���fv
�:�|�%�)!��WNYT��.E�	�I��4Gk�<#�����ȴ�u$�
[�=Ċa2��_��~87&�=.��%��{]35`h>�t:l ��8M�I0;_��i`P&����X��Ƴ��zrn�>�=}/(S�LEP�	��Px��S�D�ҐY0�ayґ�'�d3�JQ�6���|��^A��`̹�@k����3���M*q���D�Ĉ�Ære�%���H�z�_��޺�V_�ǲ�Ddr �:V�8Ī���$>_/v\+WR���|��Ľ}�ۊ,��Q��/�r���;�w2���;�W��ؼ�|K�\q�����i�E�v�=5���Y
�c0��2a�~�hS19�#�:�Q,D ��D=�D��M���k�7�s��o�P[��ѽ�W���:�ՉC�~��F��j��-�0�r�MK��{����o�1�5���̸��������ߔ�� �dpD�v�!w������'���̴�w�2QF�P�#�m��n�g ��2�O8�u^!�2d]���p��x�9�p����Ϸ��N}�V/J��bH���5,ӂ6R���Vi���%{�Uq��ͽASv�s�j�T*H�t� ^[��dh��d_pc���I�����#���cR@��$�����l?��a��:Sn�s���}0\�4��T��!�=�7�x=ֿ$��yy�̡7��i�y������Y��X3!�繖�:Xe�,�	������j��}ѕ����
A�j;tT��M�`�u )�(~0l�4�K��!H@l�&it㞞չ�<
k�}��p�K{�0o`R6߰��V�ZV 6j|�'��|����Wr4n�q{eR|�n0��x�Z�0��4�4�Yf\�
�q�m�S���IGox9�D||��vyt%�h�B�{^m/�"̝u����vy����<�K�$����]��z��24�|C4 ����	�=�Z�;��fe;�ᮁ�R���Uoj堫�*�6�p��͋Y�J�ٿH�<���өNi���37'��Z̻VIK�MH�*:*������#��m*u���Qw�u9�.Q|-���w~!΋\&ێx�ǌo��$	��r@-|+-M�&h8]�����z�Y/ E�7a��r���{�`��̰Gt|����l��D^�	��y�<�( ��\�Э�×�y��|�\�K�;T�x�#t Ӑ�R�V���1�0����q�,��֫�Z��LQ��&����k��-�6��'��E]��rip��K��"y^�ˆ�W�N�j�띊H��}yҭ���\NY{#T�˙ݽ�0Nmt�K�}]gť�� ����B��-{,2+�� ^v���<�Ro��a9�C��dr��0y;�G�G��"iՌX���b�]��\��b��kA���N谤S��B�ܼԥ����Sg�4��O\3�v��-U¯#Ϋ��OM7w|��p�3�9eT�T�tup��ٜ������A�>P�>�m���P��tuP%�_ :D��LK�蝽����7�fF7���w� 4��W���Am�ϖ	/N�:��G��ʡ�5m���>����|4ߘ��F���♰����V�K����#����+�)�K������<�Z<e�I#v��D�˰ՁsVU4_2!A9�@_�0���KB���>��1�M���ƴ�m�'�P�f1���03�����Ŷ;Az��C]�Y�|�;V(�"��:ʜbxC,�5�(�(������؂�(8�mn`^k]y�9�.��]$a�u����C{s��r�	�H ��ڔ4�-+g��%�x�+���h�
~/��c��p$2�����<��a,���C���#�7����սy�7+F�8*��� %C;�Y��a��� @�'�+<u�௏��/��REQH��ᡇ�d�����J{Օ��%�U��j��*���q-'�NԳӛy�hU�nZ�4
�)���O8�4} ������QM�QvJo�'�ģ���zěT�z#���$g�qU+�$S�7��[w&dY�u�W����ȝ1e_��&q��|{a8_�r]J�xaE-u�V�1vM��(wG����0l�W��%�	��!^V�U���`߮��b�M��ۿR�坄�Xk/���ׯA��s�����!re #ώ���p\Y�l��݁�%c��Ô5{7a�U�����4Ȋk&�v����!b,z#7���m&U6s��1������h�RL�A��<�V�iy\����D����;��_jqp���mG����~ꮮ��*�o4a>X	S��Y�?-ğk��-)r�w����9�?���"���gF���La�bm�A���m;h�T��68��\A����<y�����-�bʿ�[�$�(��@�d���ߧaq-R�Iv����]��0ΫeGƵ���:�ݲ��{Lm��ύ��WD�,�N�xѱ�X6ǯ�ئ2�tw=bB�'[�I�?���oʗ!�,É vx������z���Y�~�=�vQ�d�����n��|�_��s��X��\�d~�t��,_U����T���n�K�+ܢ�.P�+�/���Zd$z��>�>�eM�ѥ�1E�#�тl�@Ǟ7x$4@�$!�X�L�wqz,�lO��iM13��CB �˫�2Y��F������?�б���?�	�t�4�+ 4JCg�cd����x�)�K+٫�U��0�b]$���}fk��-w���	i���>��.���q=�H�=de7Qg�Z~Y٘'q^�j�ƍ]���fR�LdX�#*�S�3��w��݈�&y���t���g�?ω"H(lx����e���Syi��¢?�T������a�j^˿ἇ�:���q����)��5I~���SU�~�\�t�ǿAq�٬Y���5o��l,�ʴx;�����JZó��Q��+��^��{M��wHӿ-*?�Y˪�`�;Oif�Ċ����Ui��Q���p�M����MW<�Ba��Ŧ��3��tn��0�5����i)C�oE��_�������z�WT?�܁������?z-쪭 ��3"��Ǽ�?*��ؽK��k<��~Dg�L� a��(�s��\�۪�/��l���_.�KnbR��,I��r����*�p�-
�Z�%���4���ڤ�D�}��x�'�1�\8'�Ϟ;�|�ދI+��\�*��q��8}-14��ئy��&�$~�.���\5�j$�L�a�
�O�'�=\�=^��F>��C�ѧ&Mea�9������� ~�Hq�uK�j��/���l��`��w_A_\��ќ��HZ�?y�m'FG;˓B<��n�3�KJ�c�n�=����zu��R�w�Ƽ�naECM[o��뚊�ѥ�k� 00�ìל.�\�$bRr�d����@���7�Z��+P����O���I��Lªo�h:	r��0��Ti�,�6.-�d���AA^�X ?@R�a�������g���A���Um�z·�!fA�����辧��.�0���RG�3���<ff��ؘP*��08��lvh�>�di>����g���)-d��1x��[�ɭ cXsJ���2��Qb�1x䟮����n�!ji����n%$�"���F-<�������ǂnua�|�A���~�r�uR�뀢��E3 :}^YD�!���? �7`g7}�a>d��E;�%� ��E���m!�!�N� �V�9%����u�L��x���a:��Ji��sf�<�i/��%ܼ���D(�z>�&�X}{���T�1V' �
"8�k�Z/2�K�^�Wb��؜b�i�k+ц��W� ;�-v|�X�1���~P���T�o�=��*�|7���r0k�1�$i��0N��������~x4����P�'g�B0��By��S�4{�����8���p��3A��&�A˸y�Z����e��_��,,�Z�������eg���=s��ì����e�ˀT�
��	c���V�΀G���/�L2����(���Hp���S��3����(���������W�� M�tH��=�y�`�ʢ����ƫ�L���Flh�BV�I!Z���+�&��� q�k�:���3�x���{o�m��ԟ��\������"�o�#�R��Ŋ �1J6���_��~�MD�M�����#`6I�T0,ۅCG P����,3ha+՗���m���[�$��|@�5��Fnk�ɐ���b�r�\ȧ��rWL,�A(k��(Pl��E����'�H�N�P��eR1���x^�J��;�����$�p`� ����<����Sn��;�k`��cA��G�Q���-�n�anh\�
�c�������?Τ�za�)��&nE-�B�'�N��w��l�.����M�H�Ckߏ�@PsKŃ���#W�mn�S�����a����������~;.����_ i�zP9ɟJ63'�U�p]���j�X���)�t�AV���w�7�*�����6����8C55��ɽ%ʡy�E�R������ A�`���F�͈թ�lDq1�_~�L�Q��!���j���һo�_��OD8�b��v[�&�z�}�
��ً$�6��N����BR��yk
�bDe_Y@|u��P����B��Xկ���+�C��%K9�Dnt�uv�_������ǟ���~o��N|�.�����TN�lV��:ÁǞJ�B��x�da8��^�L眘�ocmo��s�}?F�bw#���q*�&�eth5��+�^ګAZ�\�R1����r^��
���ˠv��R��GK^�7�z�M~���E��W�Y��{8f;M���De������$��T������k��G��<ä��I[���N#�`�)�oi����e�V�x�ⴶ3��3�W9('���7�(V�o�P�����D��� [P�p�?�SQ&���#xp����{�1����o��XSx�ʾ�g4�"����՛�Jl�8����du!ئ��ք O����t�����W}��&�;�����p�c ��`=������δ`��롺F5�>�����۟�vK̸����ǒ�Y�� k%�'1�>Œ���R3����;��O�貎�ٍ[�Y�{n.^��D�V<_�8\?�>�I��%�F�wa���
{[/���� %a��T#jn��B�{.pY�p�C�^��g��<]�����Y*u| ,��ߧ�ж̘���I���(��d�]�������؄��&����qP��Z�dQ>;�ۿ�E�d���A��'��:�i����{�ÍB��ρ�5%MR�(��ld��w��uŸ�P�3�`~��꡸�-� �����~	3�ْ�\j!���u��:6�������4J�E�}B�����=��>�C�Q^4�Fk����CiyU)\c��\rŠJ�q#�z	�=�B^v)J�ߏ��1�L��~��d	G$/����~/G���j�8J�'�OI�����7���|�<��f�Оf�Xߕ�5��J�V�>�h7ALsVbZ	���_�-�Ϟ�xX!���k�'y֛X�O��٨ �w[�s�{��E���!N}�Z���u|�^sS���t��cX������2�Ե7�^Wx�pC�A�	�ڠ�(h%�|xr�}뚥�N��g��trԇ���<�Л��ߨ�A�\���b����
�`W�h���4=٤6�-!�Zaq�`i�@�?nܡgq�9�x��倜˚�;�޾��G�9�{��bbK�qp
5I����T�uV����~�O�)�B:�#�d��hV�ҒUWt$	�}gp0�b��6v��"���Z�XM~O�����+V��*�#U�����#�	��Ȭ�W���1駙���A���{57"�5`d7�55��� ^]��A4����!�?E��)�o�����5}ih fe��C�UI�C�<���Gh1��r�����]�dke�f�q�^ٕ��ʗ�k�頕�aل��x���/.���g���w�8���3�W�f|u�p�T�!ѯ�l��2z�Y�($mB��ixR4���v�M2��k�=�9�������Ō(�f�tu�I�㦑�f]�ɿ�2��/��d�
G�d��P�������"
ރ���w<oK�crh��2d��Ć-�cq6��ŏ�Řh� .Y���E��[�6�-F���E���R/��0�}��mwEz���W��?�a�}8hY-woz�U0X�W�W�۝#��-1��D���X�>���"�
�<�p�M���]��s�۽M��o�Z�Q(̒�C�Ri�TCh��4g^F�>���b�.ނ����DAQ��59���F�"����_o��VZc�·\Į��r^:��p���pkeI�Y�\����o��Ϯ"4`'섯'�r��qf'�"�^���a��^�OB�?�	���oa�����5]��Z6�q@u ����\�E%8*v_���~w���M_�
��ޏ���`�\�\-���+���U1mDh��A�I�0� ��G����{$�X-���HX���3�0�vD���m�(慾��ٸ�U�Sӭ<�]
z{�:�H�@��j*��i�j��	��@��[m���R!\`1r+��WfJ|d������΁&��P���+jK�>"zVh��6��&�yW��z��Xx �su�8�x���5h���B�Z��C�7o=��ÖqD�~t�,8�-����Lc�����\$Z���8
%���k���2�1 ��ȒA�*�̊��@�J�Q[	�X��4ш9�;������3�����Qˠ���Q4����o �v`�C��#P�O�[���7�R0��#�<�6����=?�EvY�P��\G�-Y�(&�g]����w���A��v�RjU�i$�p3%��|��,E��)�j'����H����%T|M���޶��J�7
9� �Z-P܂!!�\usC��wmt'�����L{�
Q_��x��2���b�i l�(���u�[5�bX�� K��v�cH-v\t,�(�����*C��<���Q����l�#P�,�����O_�'���n2`�%P��<���
]ß��.WJ�j�dX,�EM�]�j dT�z�ن\2�C�����:�x����N/2�����+�]��;�k��
�W� �(�y͛ڏ��^�YH�O!��E'#m�j�(w�i�9U�鼞� r�"
��.1�S{ ��b�A����Y�׫�IײȠH�NLr_�C:qq���W,e%���X����^�^�$�<XM�-�пo�]��}Ҡ�5���}�y섻,�i���p���V��9�fsH8lH��r���7��)���b��?�8S��/%�$��D߸�=?�E�{{���CM�>p_l2?<I'���t^�#U����
�I�\7rx��|xm`8^6�������(�y��8��ͷ27�Ix+�A�{WrPE!|YUC|�E<��O�M#�  �T�	ctA�d�a�|H>��\�c_3̅6�cZ2����d]���� M��v~`@�@�)�apZ8�`2�ѕTq4�g��cH�p��a���1Pk��c�A�NR�d���&��V�C�f�՚�Í+sSa���HY�γL8h �q9IE�hw��0)<G'�����������x����H=��J9��o��-�'���'ab��k�*�*{)�># XFD��VY	p[`�V:ܾ��v��Uj�5&����ZL'	66&��NS�~�1[HB����gQSS�+�*9�(�+�3�@�M�;u�t�X�Z��m�h}:��r��7��:��:��4��7�	v�hS�j{��鷈b�S�-���:4���rG�e�ʶ![�	��`�<��A����}���$ڥM\���?��D���s���,'�sΪ�IT.�'��)0�h<��1�������3H|�R�M�V�b(el�2ױ��I��2A�8�f�CBR�i���^�:"J��N���{��������j�Q��L���=Lq���t٦��zO�eq�6�9l4�A���<zS����8te��+�����>���@Jb6Ǘ�i0�?d��iOI��N%�
�5���}�h�����=O6�zFQ�h��r��s�w(P�R4"Ғ�DGt�������_��e���j�z��
z�I�)#f�� �_��#ص�PL	��Y�LH��|�mf�v� U�r@����N�Q,C���p��?֗�w�8�θ��_��C�Q�FWb^�/p��2T��(n�`K���u�EB./���*�	�G��qM 6�I�yӼ�L�|�T���^߹�������C����ݜ���a���2�(il~ʈ�w.�EtP甚�� �w�2����4�L���*a����:�e���6�LF݌���4�{�D���T�x�#Cm@�v��/G<�����Z�9�u޴�C�&Q7��&C_�������B����Bs���E�����0��L<ӊ��W���e� ���غ���Q�+Cx���Vr���N�+��7�-a�������Q��O�Y�TVaI*���?�ߎS�+�`<�	�B�s�z��(��V6t��r�w����ͺ�D��kfp(�:�U�=qJ���9Y4��kX���9Q���CR΢:c=���5Ҷ���Qu�E+`�0����R�P�`fIz�=n�a�����L��G!2#����n���P-�*ҙ�B��JM�b����>��o@�&W�+�=]�_vh�1�Cyиc�带CL�d��ͦ�t�x�e ��HV˘,P�<<��Ѩ��E 
� N�¼ό�v��; ������F&�
��)� _��ϗ-p�qT���Н�T;�/�?e)o;�4�.��}f�Lǥ�=�(�q�bY����7��l�S���S����/��}�?��)���ކ���n;k�/�ι�\�5g�.|H�#y�oz?��k�S�+���qE����(~�'�`_�!�p���ڢ�)z��bM�d�R6�mX&�%�}������	Kr��w�	_F�#/+P��[s�iL��KLU��A�U�����ǀX��@���Q@��z6��I���q�m�q2N�����QҀ&�:V�E�%��!(���Y�{���0���o�7�D��ĭ'�(`Z2v��t���CN�{{�+�[�z���lIIx���SEF$�zć��N��)��\����Uz-��},3OK�����ڝ���~Y���*i�xJ�ף�g~���}�r\Iw�5���c�_,b��H�%� �x�z��V�/O͘���.$�����wWc>�ZKi�k���g���c��
�A���>"��L��ol!Pdq������*D	����)h6�;��_*.�<vj���e��X�6��g��׵J���V�Kn�aVb��)R[��H��"8��r��_�aC���ll0M/L�(P!`4͕D~@Z�����Cm���HJ뭒��P�4��*]���(U��9Pe�����/��Wr�$�ԉK���XI������+o���.����ek������y��w�O�O�[�mN�0�͓|ܳ��d��f�5�� ?����<ȧ|��Hٽ�Mܢ�:��>O��0:�k���	k����k%r�����?V��Po��
��u�z�I+��� ʃ&ϣ��O1_��j}�o�H҆��;a���[0ۻ4�T�������_���ѓb"|��3�1pD��=X��?�M|�+�����#������0�K�/���dF�ג�Q��"��Sc:Cc��/�T��_�Z�� ���5���# [D����F�$}�#x�?���N�8d�(�P�C$rPIҳ�BW�ܭ��a���OQ��)d�(z�.9}�)hLq-0��>���br\u�MgWs�7�W�T��_�����BAz�#�����9ͨF��̓3;0ν�':V��dUt�� ���V�����\/Ls�u��g��?{�,ڥ���|_��c���H(��:^2���+��92�H�+��Ӱ���ǧ-���<���b����YQ��7s?z\��a]w�N�َh~\�1�_�Ӈ�P�@O��BL��>��w����|���nf�WH�{[.;ZM��0�-�t��?�{�8H.y�I�J��$��K��"*�)>��oU��.%ck�Tz��7���.�g��We�GV;�x� "X�j�b��s����V�b��m�ѧS~`'�-v�rp�#Rr��ω�V�L���l����Z��� Y��nN��g*ȴ6l[�=m߲�- ��|�R��Tk��a�5o�2\�����ǷS��!��B���`��ަsO&$�bԺ���(���Aͥ�i�Ye�+j�I��ۑ����ӯ�˻���)^��?@���ۭ�ր������}Tҕ����/�D�􏮟��#�M7�@�"<	�v�6��;UNa�v��0�ѥ~��+۹Z�v�t�)�o
"n�m��T-y�`�|��W����,��UZqg:6E�
����9�d:����Q��p#oP͑�@"���SE+Z;���ID)Q���L[��ov��>5�x�{��l- +��_- >h<{�0��^��+N>����@8<����+��jb�X�{0���P���o���у������� ª� _�F�z	bT&NJ���Hvʘ]k�3���� ]�V���K�6ط�5��H����Mv�=��w�D
�
˸|#�jb������*v�d2���*M:9$Ku+�)׊NK���0"<��Djx6�E�u��/R����Ϫ�UV��HA��-C'3�
�AYU1AGrX���R�8�&<�)��.��3rE���pT�{X~��`J���z#";!��3Y��(��78A&S��sJ�8���Kv���h���d�I���;�E[���B�ם�������K�S���l�K��Ōc����n�/�0�O����EyPB����IO��j�ȟ$�� �@\�b��~�]�iy�v4��s�5gX�e��O�����j�J��S��{^P����Č~/P�*�d|}[���Ʉ���Mw��`��5�/����nο_C������Er�*w8PP�W.������)7L
�8�Ế�~#�9��nsLB��|��q��_EK��^ք�>��K�õ�i�s�+E0e�D�eo�M���z�P�����!ſ�vGݶ�a���M��\�,ȷ5��"�N&�b����<:9d��C0���T��I�!��5���u$�֦��h�gu޷!A��рˋFr�@j��t���LCh5� J�mu�݀��sp�#�ǣI<��Y�;��7	�vO��tI�pw:b�r��B݂�ћ5
A]ci��*�ʰ^���g�ЄC#Md<pT�jA�����+7��*9���Ӝ�l���g���j�h�$Uc�� ����$�_8G�3�"JN�D�����I�?��o:�+f���6!z����8�e�V��B��h��%9��v۷�w�q)�̯���"!S�f��U����y[F�4u�?��qO�T.�W�GC�~�
�BB��"G��!�M�>�:�~r�B�Kle�B"xG�����dY�d��NǺtmS �I�s��l	E���U�Xq�}�� ��N��#HA�Cm*�IA�PI�^��g���?|��Bag�Y'Q<S$F�(+���t�E�f��Fټu`|�!����#�����F�ݺ���i�M��յ���e����+��G?ZltZ����+i=|z��[/�b#�Up"����>�ՌbV��~�=�b�puϗI ��x�9�i������'�ar�چ�'ys���|�_�QN�����yGb�(�I �̊��kA�������7��x-�%���Q��m�(+�C�_|����6�0�v����Ńb$DQg�,H&��'�#��;��I�d�[�!a���v��/d���r��E+��^�D��6hke`_��}�39&�p�q8��|�q��xMz m��kx�I���|ߓ�k�TLg��&ԾK�lUD/�@a����ϵ�]}���L�
`H�ST#�l�-��P_�z�������H�n:�d��F_&k����9����w�L�C��^-�kM�5Õ�/���1i�=�Vp.�
Y�.���)��q�F��b��o=�r���p�4��f��cg��뉔��ZY5�K�#���P�YbM���T)���aLJ�	\Q(�\���#V�W�&�b����:���.�eϴU�~21rO���%rI�u(�7 �5��%M���1�@l���DӢ4���)��8�(�l�1��۷���p���c�1�R�m��<�3����[�ٰxͮ���r����cY������\��8�m
�>��]z�g��Q5�ZP�Q��q]�"WRR�V����#�x;��v���B?�C�ZK�q/���a���;N���#a���m��^0|L�+Q�ܪ�ut��w�����a+:��p��K&Z��Ȅ`m%,Q�hS8�Geu)u-���K�`���QQm��I�jFs���F�@L׉_�Y�� ���1�=#ߥ�\3�ڡ�����d�8�0&]3�2����`g�R\��>
126�<������ %ʚ�Qn|p5�ȵ3�:M�gzP�ǁB�i���2�����QlҮܷ��M0�䪇^�ڸ���ddXA}�@(���RMKy�-�S8=�ܶ���I^��ec��X�ޘ�]P&����>�So�eX�yr���UHcW-Q��v[k�B������o�E\8�N4MU{��[OApj�'
�����F�+��Ӽd0�k��ֹ�́55�J�*����QrJ�݀μ��,wy���-��
�1k�.w�Sl2I�iͮ��)�zY�A�ɭ$.g V��[�������b���[����c���tt�X�׮/�[�6�Պ�=�͕��	Py�ӂ���^��ר|�U#��������1�!]����8�>ˠJ~��"^a�yB҂�t�wpC�?����4�`�ڂP4�I~s�͓��U����<����vOg����i���1�������L� �%��a jo�fDV
6��y<ѻ���B�.�5����������Mi&@����h���y{Q�;�V�]�l}�AC$N!���iO�����k�}6�U�3ʎ�鵲-�C�J��:}K����y�C�	Y�,�Si�Q޵�?��
�Ƴі�Д����G�^,����H6AP�kd��J��wo.�"�5�Ԕ����3�^} R@�����o d�یg��aκ\ d���!�&�ŗ��(
��H�/r�W���׶Q�tb��U��C����pQ P�kN�v߇��P�+�lή����h��)��U<��!�Ϛ�҆��+xÑ�5�$�ȉd���੦?��Q流}����8�sz��#t��s)���`
��(X�k�累1�ئ�ݢ����_7lq�ᐳ@���#�r��P��=~��k���MHoyS���S�QE�>{D���&K����[x�����A&�i�>�~f�a4j�FC��ӽ�cd}}jv�s8�E��@�O�w�L��NSd���K�v����
s2�9�@$�X���}����B��"a~���H�s�{�:�8�cX�,o/b�\�L'O�jh�m�Z�!� �}_�ķt�JM���I��bZ���u�%�6$����l�!C�!I���m���O����?�^F6c����W�:-�P�ع��s=�qd��"����.��gpo��C@���ۊ���j��@$-��'h9��_y����H=��~ w^P/�4���D�=6cH��QV��^Aج8�-�N�;L�����}�)d �ZO=��İ��	�kDHՅ:
H><�g��ߥb������W�}"HO�`����D���l�.�L¥H泌�+0�JZXF%u�|�����`&��}6D�JL�� 9��<ԲHŊN��r��Kc���ཎ
���}`�0))U�сNhAC*�!z�Mx�度�P�����[�e+��a�8��j^��ӀZ4:���X/��8("	Gϥ����S6��7m�bS.��)Y�Ge�}���^�'��P ��%q���X��f��������CJqR'!ZF��,���y��dI����;�5��Ӏj)�In7�����%a�]Ń�r�W���x�������gHyh�>[Ӥ\��K�K��y��[����I�q3�E0]��d�p}!�M�@1H��w�=z:9�0�)^#�h��iݬ�M<|R�J2�E�Mz֕oS�P���Jع(����-P��+'��!0�OE�����;�OXNü4��n`<G!�,���Y��w�[�蛑yZCN��l�F:��#��˓����Q�t����#�W��b���$�K��ţ�o�׺�LWM��.=6�b
�τ�������ML7�b�_/4_�mch�;�&�r�-4 �-�(�e�{A���oX0�����m�^	�^�j�OAѥ�j�;8{��*)b�=O�h�GnP/#A/��"s��WH`�N�:e�K�����U��ѣ�WP�~�z��ąk��+ظ������N�A.�$#�k,Wˑ����&��ؗ�1Ռ͊��,+�z�Y�4)�2^wa"�e[�Mf���#�F�ۈ㷬�q��vMA�|�Cp��咬M�LXEb���I
��^6�BɭK%n�l�y�H6�:LČ��/���D[����1	ȅ����9�C�X����Dő���v'��Hk *jn�-�� ���Kψ���Z�fR���<,s@j:X�é<�o	5������;��8����+"� �$��ېh���&~2�`��V���-���{ho�ү��6�5�	sՖ_�4P���?)�$b�3�ڠ9�[�I5ʯ��K��f8ь�Yk&[Kq���#�_n9��F}���8��$�t�w�|4X)c�PuH˛����r
�c+$g�����
xO��:�觔�u��I�OM����*Զ�܋<y��Ldm�Il�㥦�wW��>�'��m�3�E�MA�)���1��4D�dA?d�K����Ȏ:�ж��Ua�	�������0J�)msi/����z����"X9�������3&�'O��AX�rV�Zt5Um	n5����ʯd]0��^�wU ���P�mU��5�`�P�Y�Jd��:t	9Q�� #e	,ܢؔ��"1���.I)��q�!" XG�a79����ixeH�Ù�*������Yo��Q��l�UM=d|u������s��A�ͣ-�GX݉�]<�7r3El��R嫰��p�?��r��Υ �ݞ9(�-A�݉�}��c	Y���
���l��̌�'\0PN�n��`":��=�M�'" �Vx�] lo���4�\��y紋|F�b�*SZ��-��v�
)����u�G�BY��Ϝ��~�1��fl+҇wG��@�P��(f9�4x���B��ֱ��US�����IN3�k#�U_��h%����z|��>g}s���4lL���2��[f�.�`/uC�����R��خ�K�;������O>�K����0�+6�!F��3tHy���^r��n�#�Z��C�`���&��՟th���&�D�}�w���W��GV�=��lƏ��:��X�[�7Z��@�{�8]��ۦ*y=�K��� 4�\ͩ��͘o���,�Y>h��0=���&d���z�(�BP�R�v���Aҟ5�d0�W8�R�mxOu�!E��v2�1e���c4�,���E~ZөK��?�>���%klp�Wۛ�ժk=Cܗ�QM�gt�߅-�^���F[��)�r�4JWF��f� X��Cv!��{��t0���Nh�Ȏ:��P��%v�D�*W*B^�]jF^`d���?WC�"L�դ�%$��܋�>K%88���Ʊ 9����!ƫ:쌍wb�?��A�g3S:�Q�H��"�MG�����J4XEz��j�o�#�����P`�Eǘv����a�/�
�w�pq�|KN��׻2dK���R"����2��ըFf~��C*)�-..F��k�#*��D��[C˰���UވLV�S'��p�ʬ��E�n�h�+��.P��Pso�G|�^�d[X��I�����ds"������!X�G�?���e+� �9��l�;���)xb�X�{�=H����h-���U����y� �#e�?QY&��ʏ������aߺ���H�C�hY�
	YH�����IJ���H9�i����@k`!��6k7�o0��M(E��b�r��Qó5O^���A�]��#�'�AA��_��@jA�A�W�.�Q�����\��9<�%�AYW����Ç#FME��u6L~�>^W,�H����>����Ei��TR�@��ֲ9ys�g��{�j1r�3�]ǵ¼�4�c��K����wܟ�����+T~m�/�R1)+�OVC�C]iY�v�B�U#֕Z���⤩��K�����r	�]�۹~V��0)�k��<�	�-�c(��¨��1K�6�,L�hd��Im��+�D���T
�ǈ��؆�9�]L�˖<Z/��-��L��M!ؓ��}G�,�"~��2�a�=�ya-Q9��Q���E��*&�t��w	H��?�w�Sc����2²�5n�z_��؈��ŏH��\���E�I��"Ƥ����ll����ۉ16z��`��4ګ�T/�w��	�P���8�n�e�2��P�X�ǻ��X�Ha�}8ܫո,)��j��7��]�z��E�(���A(e��́�����,cj��$��e��9�S�m/�V�KU�J���Q� |��i��3~�oןv�fH��s�����é�̵�
ީ�}��-�0�XZ0,:s���+(eM����:S=`������f�B+��Bs����!W������8���B.��H�����VZp�7W�;���]���Vb�
R����8��s�P��9��}�6��n��>!Ô!<�J�4�d8޾K�1`{IƐ��JJj1s���X��\E0y� :LW�������lE��.���0��Q���|oo*)?oƻ�c0hW֚��l���	{e ��p�,	��~噩֏�g�聝��\9ի�d+���b�='m]�h�{��	?�4_,���ir�?@(��/8�؄��<��˼�*�4x�02=�jY����Y�'5ʐ���j/d��"�d�Y/�wd�g;��#<���i�-|�^B��v��q��k  yְ;��ԣ_@�4�3^��_��$AV^���nV}?M/�S	��EAI� ���"�?������?	�je�l��$��lFn3��\RЪ��+�߹;�Y��8�n���Ou31��Qp�	f��%�QV�wBw.(���M��4���-Z�A|�PtuޢU��m�0i�S(�򄫦/����|GlQ���-N��a�'�5�]Zh���z�*��X�$)#�)w��g��k��FaNm4z��6cX��r���'��"�L{s��)'OýߙΦB�jr/=Nw�+���=k�}��O/ݫ��;�)@������F91B�I���?E��wĹPV���!�`�Pz��,ڄ�{ȼx~���v{�v֯.�\���(Bx�CU����b�}/��4iE�,��.|��j}u��0�_�:$��F�@�}u���l~4wU�Ed�
�����2�k���f���^�����|��Ԅ�]�bܼNH�?`wa�e�䇆�];م ����,����͚j�I�0��XS��(��x��]?�ѵ#�C�T��_Ϩ(�d(~�����J����~y�H����m����!�V��$��)�w���u�L�3`�v<;�Na+�v�XU�=me/����?����g��A�9��O�2�b�'�ʇ���ʧ����VӅr�b86���H�;��2ư��?��._�J�`k�����F'�����%� ep��_�d�[(js�ay̯p��n �˥$ŅYa��f��І
��t�
 '$�_���8a��m��������m 3[Dwܯ�|�-�c�-w��G�H� �p�Qry�!���~x�%no� i%87�ލ��V��A��t��v��IN�ُI�6Qa���2��0186	,3�J3:2>��-^ �w�s�iXa��}���� L�{-vwȶE���e_s2{��!�0*&���8�f���=�X���e�o䋅L��zĿ�މoI?/�B�Qw�w�=�B�A��r���7����+�^SwX�۵8�S6���T�I��Dצ�4�_����M��|_�,fRp���%i�����r2m��(6��8�6ֳD3����;�D�!�`L�j�Dƹd����0��?0B"]���	��a�B	C]_�Ҩ����V����^
��Huk�����vϞ����;���] ��+�=�@��0|�S�
��<�N&��ߌD�j��1Jn�ZL���[��W�3b����X�w��:)�|Je����\�?I8��\AN�孊o�Tt:��?Z43�x!��(U��'[��lD?��S
1�V�2�Lm��P	]��D�w�7�xc�NL��)�V�lC�������輾q�Ə<،�Q��ͷ��2�]g#w�o�dj�s������E�����Y����I���y^3�/I�8����u~����~[��s��\����,��<ʪ���r(WS�iT��-�&� ��ÉH��[q3�I��=�ྡd�ȚI�U��*7Ԥ�C�\�����d>�C]���;�g�@!���`�_4��:���O�a׏���Wh�7��:_�ؾ-��@P�{Z�QԷ7��ҕ{FX��K��#x��̨�t�>�"X�XCD���Ml�@��r�c\��K�v"+����E��P�j
e�4����S�)<�*����W���V����*�&%�4��w(�'z ��|?r�_$i��1:5[�`gk5@q}]�$qk`��\���a�WWoK���P굩�Fߣ *�����v�~�lư�sFf�{��h�#/ �xۜ
������w�|�����A= �L�;�6���W�kv��+x��~)���^�y�N�ڵ�*�d)(��ejx--~�:Rreߔ�S�
�6�Ԗa'�L����1Q5]�Ɣ�?���D�y���!ЪY�S�`Q���@v�E%�Ӳ�F�A�_{7��8�18%��:�P
i%�Ά��n���~V�Y�E�C�����m����g��o��Oc��[�J��|�� �	-�?2���KX�E���"WaD��l�^H��]��+�J�آ�Y���׮�z�DDB]w�gˋ(��G��������~Δ@Y��U��q���kՔBZ�i�w�8<C�j�Ȏ���IҶ�M$�c,���׍�Yo�Α)���k��]���\;9���n�K�@���9��2N�m@p˻���oP��d�a� �'m�g��`�쪇�P9E3e=[:�w��K^тk��	�Q�|c�f�t;���	)2ÿ��3q��uu5���Aόcl{0��jE�A��W� X���d�=���Ndb����E-G��RI���A,��^�lR�-	����Qd�Hu��pun�O��$�)��T�6g�2X����ukH����`��wN6������$I~NI:����������C�!���š6�����"�wg�W ]�Q�RO�1j��:�	�����KL�b�^�[�d���N�S���l҄✕;�F�5ny4���z���>�'�z_�r�Rȼ(pm.�|�i����_1�:�݂�I �)9��a��M2<?>�-��������|KVV���!�(ײW����a��-����j7��cq�W��h��4�JJe���*�_3���g����`�Ot`��#��F��1ԑ�J�yјv��־UX��b����t4��*M��3in��W4��T�o���4˻dF'gA7Ȋ ������֜xV�̼fLϏ&૬��P[��g^�y�^PI���պ��GU"I+ �8D���  z,��T���|�5��喖��D�I����"���P�7���ot�76�|�����Y�����CdiW �LN���g%rc����d��$����B� ����#԰r�Vu8/�CE� ��{�+%�L�����M�(���_��ܤf�r�!�
��X>�D���ۚx�t��m~�hM,]Iz/�	�#Y� �Ϩ��]��N��Jh���\�1�°�Ƭ��� E�#r)V��*b�����'��;
���)�I��ҝ�i��n��%�ӱ=�p�w����^��b��ؠ���-]�@
��ٝ��J_��Œɱ�.��T��Ŝ���0�?
�}��X��\}�� k@y�oWƅ�Q]#4�slŦ����B����E*�f��~B�¡��g4]�H����[pM��ze`oc��[��	�l��lQ�X�s
~�g_aj MV���r]�����؆ ��L���$�ة�l�(��~
���0M�unfxi���Sڻ_�ƭl�&^R
̟�_;���kX{�E��ÉG�r1wI�<�y�TZ\M^�d�5*�X�M�
��笿�ᙋ����ڶC��W��|���B;�W�4{?��#�Ǥ?��]��X:|C��{�K�eο6u.R�����r4Ùe�r�z}�V�-F����qŀM��MT���ڌ�q[�3�4����a+L!����=�V����F7R��6ͬS(�������L�*庎ό}�n�P�@���8J(���u��&/#�>@�%G��Z��-()|�ˏg��k�d��":���6�*�T�}'$����K�v�-�ل+C�=�,De}���jY�ں�I�^`+�G�TZ.. DO@9JO5�: W@��P��>]��B�6�����U��A�(���2k1����dCqNl�%hv�1�A-#�4{�2T�z�x��	K
���!I 2��[z)�'���J&����h7���x��"��uG/}����O륿W-{~%�����+qbB��Jb_�O�^b܈sܻ�0=����Ǧ�)������2��}/����M��
r���2���;�M9ڝ�����S��0�zR�=���ԙ�4w�p^����R4��(`�8^7=�1�SG��0��D5��Oxo,�e�K�V����]��?ƅ�����
�JIɘe�{����zݗ�2N=�G-auWQ������]���^l�G��}{�$���*��/��kç�֓��t9I!K0X�B%��/���Y��9rS��nt�pN��T[�ev��$S�����`�}wZ������i�$|���/�y���Y"ـ�'>"!Oi���R�/�).�:ԫ�,����{��v��� ̿X^ꂧ�l,[��:�F@}��/N]�EK�XG�Z$�\rm?A ��{�)&h��^,c�:����c��<P��^H�!�αR�l�ۃV1 � �I8�n�Hҳ��K[�w����+��(�{��8�\n�����2/=Нiu�Uj��+�$K���B��g�BN�_���V�?��b�sħH�͵����z�\Z��'��l���f�$���: ����3.�Y_�c�]ú��e�6b�,axVy�+�C̚,���vJ��u�����Ӏ�U�h.w���k��;�s�	��=��[s�!�b��\V�	Y���恝�?}�!�+�� ��e*=_���ɓ"�	'��BD,�����ͨ-���ޛ��& ~t'y�=��7�@=VN|��BY�)���i��8��@�1���K-����?��k3��I�[��R ďҘ�lpP��,��[FG�R=l�}%>�������-���9C �V�=\،�n�3-�.���,�9�i�?����Q�mD�?��0�r�Д���9DiU-ݿ�ʅ�L�t��UFJ��b�i6}l<z[��;�����܁��]F�~����× � &y�� �Bz�&Qo�\��h��c�IG�I�z��:!�'�V�w�Sh�7����p�Ɂdd-�-b$,J_��\�z��J��K�����fE>�M���1Vl	�U=v�Cb� .�>U�9Q�|�oY�G���Y����U�����1G`�H�u�P�?�g���hV���F�	a������ڍ�C�����8�]�["t�Kl��BHj�MVs��=h&���w�ܥ��+ؽD �J����=oB�-�&T񒙢���҉�e�H�����K͛Mm8�q�&|0OuΧu�,T�,����P��Hr�����!~y)��>���k9ؿ9��7�b8�(v�"�Է7�`��ܬ���Џ�<V$�uÆ����0�6����K�4���Y�Ŀ��*�����ï�{o+��_�Y�!�${�d�YG_K���B����i{��B�Z�xQ+r߆n�Ⱥ�_�]���m��O���i��o�`��	>�Z7��3+(�6a�+��h�9���f�N�~D9����yq߹bk"<yOY�w����zС��p��o���e ���&�~���|�rm��V�)[o�����T�����cNf�A���e��L�����D��)��7��Z�P�ͪ�Y��q�wB�5���?��U���"���ʻ �[��7+Bo�!^jxg��8������Ms��Zoz|�4l����zB��_����'�gz�|��R����S��q���>�hA|��� �46���Fƍ7�}"���1�j�h!���!~́f:�A�	 O�nPh9��Y:�Tn�Wѕ ٪�e`W����F��by���2a(+�Þy�u�֔�.0��"���n���
�CMw�\=��|�0xb�W�r�e���P�j�	(V�.	00�E __A���O�o �]�����PFA	 �a�G>���+�ݯD�&CBC�%GX�P�j��o���\Bګ�m�B�vlU��ʺ���w�G�*�_���6j���M�)z��=c8�ٔ�c���
���sVRՊ6�`�xA�>D�
{�:�[!>|���!I�W��ޔ�n�����x�5�IA�j:��v�����l�+L:��;S����
۽3�!�j��*���}u�_��4Hr��;���۩�����C�"�ҏ`�ޞO�5��.�|��T0�˰ϐ�%h6W����R�A��d��M5ڥ��HZטE�K�?Lu8���LҚw_�Bb���oA�������h��o�fٌ�D���h<�5�"	z��Y����ⲵPC7�<�P#p_|�w�J�P	�5�����oMYqm�x)u3�{�'w��=W���ǣ�����Z���I�0�lO�5��:M^�^�>�+,�&�X������`^ �V�{~����!��� ���қ�7f���rI'����;�2���X-�q-A�+�bh�v=����R���x�.�gUٻ�@�@���A�e[�6�6�K�w�����-�'zF�`�Yy���q��1����������RI�TV��~-O��3I�T�Q���^�#��A+�oD�2�md$��
�'��\E��W�of��Lm�E[���Y�W*����	s1,��7;�$�F��R�qʢ��C2�0f)��D2�|A�>�ss��S�5�g�A���w�{ߢ�e�� �!��8;���Ƣ�l@ʟ��4Wƥ��R`[ .;٪ĬN
R7��u�͔��gι�V��|=�>�~e�[E���Op"=��f8��
�����;�*|�	�{����N�b�Ϳ��v�Y���=u%n�؋�˒�"�� }��ć�۬�XE�1�}�a��|���d��%�)+����:"S?]-�E���������m?7-�OS�:���Y�F��n�;���b�>�$�/XZ�,KM-I�
_���N�`��3qj�.4i]��bd��ӭ8C��\t�Pl��>O��
��ݶG�/��jl�����2�_�k �K�ր���V�-TO��v$ƣE�r�B���1��P��/�.�v�ڭ��	��$�:���`�7%!��[i�P!���;p�BC��3���a�#E��e��^�k�p�N�Ek��a2��{e��ERm��~
 z��ڧ%����ux�Qyү��f��6
j�����l����2�֌2e1��xP��S*'����8p$�{�ex<���a�ܘ�'w���*�D���T�?-�1�Gwr&����L���e��@���A_���$)�Fc^M�x�4ke��9��]Mc[�?~��i^
kL#}�`-%���aX�U 9�١�U��rEiN�Ĳ�J��"��X�-�X�<2m �w+�7�6eAg
�0745@��1?0������ۘ�(�k��Y��L��Z�v��t��"�ۙ��4b���k@��ĢG� �7�~��Y	~AZ;��?t����6��>.pƽ�Z3��_��9&*EV?�����=.��I�80w���F�� ��)�·q7~ ���uvg~����U*Ƌg7o'+_�"�
4ڳ
��C���%��*eD�!R��������7C`!��><��R |-U�>N�-o�!�7�kU8��U��^ȹ"D��ٔ�������4����-�{"؞�5D��j�`�y�{�͝i�T "�L�3Ew�h���L�}x��z@�ҔK6���8�q��ș<e'�t�e����2 �;h�,O�l�����9Q��kX��VH��Q�ͅBe6� �JLȖ����\�ȕl �Ӛ�gY���k��R��Of�N�;��6��@��qb;s�ˋ��	�6�5����Ef����m�R"����8%>M_���j|�6�?8��*�UI`IM}QH�F<"}��Qk�\��u1Pt 8��P���.��%dت꫖��=��g���O�N�)o��OR�C��&��0aXK�:U>�]�Y�\���z�at)J���FO��&�i4y� 0���C߯�݁@�'~�k1.÷Dz��g/�TC�$���Z`�nw<�R��P�����4/Yc�aNUx��R	.^��^UzQ�(Տ�H��]D�2ܝ�٨p�{Z4�"ܜ�}���]�!C�p�3X!.ĉ=Zjh�,6�߯_4Z�C���؍�xы$o�	(L'�,mF���,ـ�'qb}R��=���3�R�L�G�{���j:�0\`P����/�0�9�@Vi�7�r����R0���̳�jy�o&�bO�7Q��Rm�7���/�͚=���$�O�F�6�����V����E!������ٞ��a)��[3�Go=�~���8Q6Ҏ�M;�7[C�#�u���<�q�1%?^��)t�=���՛����-o"G�ݥ�?H\͑��.*x7�-���m)�$�^"�LD~ߘ�z�O�=2ٖb��u#��nu�	���j�̬2�D�yjN�F1�@[:�o>�I��_���sPJUް<*n��%Y�w3���&%,|���6��"������u�씩���C��6/G����Np�#=M�<����O�--�!�5$�j��6H��ϕ��66���9c�Q��7X?iI�Z�s�.��j���P�";(){�$��s]��rX$����4�b�G���S!�^�[�f�q��"wCy� '�����OH4�����#�frlr���L��#�r�P��$_��D��=�@�ͨק�F�GIҀB]韆4c�V�C��F88��[M)�¥�S2R%��s�G�B��>E�OcX�|�����+�9e*��!4�?P�E�iVI����o5ݚ�g:��1{1�VW7 �OD��[�Kp_
k��mO.T�3T��s���>ְaqV�~�HL�}����D�Xj:��T�IT���`�#�A�"S�7�`�c1o���8�:���$���M��߁�}tљ��T�.���B���.�k[�Kf���$�=�:��ّ��D#�֠��;� m�Ѻ]�>XiE�J}a���;h-74�i�P��M���h��@��{�Ѐn�f����V��:i�O:h*���Zb``��zCqr�P��$UDKˉV���w���z�T�`�"쿩&r��$�P_>�&n�b7��X(w
H����|Hx�H�8I^~)�Eݠ �=���E�Dk��<����79�K!{�t��'�3�y�{��![Cj�G4f	abҜRX�ٶ���efS��J� ���$����6E��2tU��֗!�D^q��=�7�����=���^�-U^n���㇡E���Ԭ.z	�=�/����j�[��=����F�NӾ�������'��6��V�Fz���2?�׾5�=���("��#i�NfnM"��.~��S<	2�E�䝑��g�
ط@N�Ʈ��H��SA3$֬�L3�� �N[�v���f("y0s!k��!Hݘ������q��'�s����=���`YU.��[�R�%~����'#D���Ɍf�ȭ�!wBB�4���Y�U���<2,�Ҝ&�/����O�#�%DY�]4[kGqYf��9t��!�oS�f�}/W�OI��B�Hh94i��璨sp7��a���C+�@L�z��Gލ��Ý��!(ӦR���� ��-y����a������� �*�J	bL�O�*&6T� 47PƐ��e���q��maH�KXWǙet��� �ʭ�[;{�_��e�Ž_M:h��[j�tX��C��n��,����Ս��5�U�Z���*ƕ��V�i��zo�%C� Ї�2d4|�+�_�7(�}��}�1����Z��`�y��<%�G�ۆ����g(���:�M�3��D��	�2��ʹp���;�Y4?*��R���SϬ:�:'a�Q���J)������D�<FC1�n�,���g��O;���ME+���MC�S۸+�5���33�ߠ˴*�Z]���rl�o#bgp�r�(�� �� �Fb��O�.ޡW�_:�6+ҭa�KV$P��'1����'^�qٷړL����g(��u;-�з�ġSI�En�V(��%���!���(�$���$�����&���c�<��m`ێ�T�!�2wU�{+ג ௅h80.?[�[	f6&�XK/pb8s�,sIx�D��@�ϝ1�L����to���qL����O�{wm����:o�~z�{��^�.�GW��MٻHw�&)g�WG���|)p+|�ܕ}�Y�c�H�7'�V\Ma�����u�G���i"�)�˜8[h�HM����ơTb��-?�,�^b���D��\�=�d�_j�bC&�;�Ɇ|��k>㋪_)��K�H�$����
2H=�)���U�#bP���0�_�0�G����V��揮�<%�\� �'q��	��/$9_#9��@Y��EAڛ��bo�{E�)�ß` �}��:m����r����sV��%<�� ��L {ؽ)ܨv��!�\�	=�J�2�w�S�v��2a6ӑ��<f�V+&(P��\:�a�ɓ
���%:����}.�������DRU0��˱4��S�B��|�Ȯ\І#���:L����KC�>�3l���L�t=���̻�ɹ^dI����[���#�u�>�,ƦD[�-%�礛������V��^�vX$��
�h�(+�?b��dX��?�-8.��I�e��\3��+����+.� �ɭs��5����(��@�ݶ[*��=~j���ޏ������b~$����s�<��K��=u0+���)�G��A0V#뭐ՠx��n��5��5r桻�j���&�,����O������&�����1DҺb���bX{�@<�9���d4@�7��Q��� ����AX`AW�Q�:�O�=�Ϧr�fn�f�Ҏ����u�C���A�ܶ��9�KF�-L�K�?��\,�_>�G�D"o��l���P�Z�tA�(`E{��b�bT/�� �HI�n�-�O�ݔ�Y	�}���}�m���!k�eo�W���2�� ZT��3��5�Rh�`���.�a�{�B&*����U	<9����t`vx�;%fƏ�C���O�c�毪��S�(h��B�l�'b{|�>���v̓�@���i�hP����2p)t85�
:My�,M������6՝,&�%��3�>%˱��N����͊!�����c��"Tb�}XN!����m��+@����e`���*T�D,�,��L�mhTQc�����c^`&���k����<�x�@I��8G�qFe*(�$�����1$rVr�Q�cUB��ݍ$�\_=���.<zN�!��qEcX����'\}���)�X
�����Iٛq�P�
��/zA����Y�`
Q��iHھ!����bz6|,�ư����m�)�+z���!h���\e�����J��G�c�JF�B�x� �����t��E-�w�h;C�XI��.��G��o#P*�sP)�U�$9�d���Ɉ�������U�־Km��Q�)��t�j��>�`�W��"r[�=�QK��N��һfC./AZ�|�B����� �B�'������^�����bT�v34U���;��b7��G�{>
�a!��Ƈ��g��UnXu3&� �2҉����n�e'���PBn��& |F��'��G�$1��izn��e$���+�|[�므����BsJ}�"̛M���mވ�1�=�+ ��8 ��l�R��`�O���{�7$�v,�m���}�tjY��w,ړ;,J���M�O�m��衁���Y�[��|���lz�ʘ!��KT3�"�\(�C��zއ���uW�B�>��NP�E��=���"0���b�)�ʱcz}� �-t����ڡ��2���qͧ�!����;�_)'֡ň2���3�QqK7�����Y/���m�ޕ��z5A�2���JE�aģ�^C81��|�B���-=�����/����4'`��1��x )�c�8�����������y��p\��t����/�X��7�ǃ��J��tlS[�����li3�����t���76�H+<��� �OU�)$)*d�޸�xo�X{�1�G45g��J��"SL�E\��6$�񗌛i����A!{��}������ˁ�R��#%�d��\�,��N$.s���{q~j\B3O WqJ�z�8�<���W��_]L)m8M�P_���F��hd"���)���[B��=��~���!�N��7�xQ�m��U;e-`��!��W��[ֽ�"��-�.���a��n&���tW5&���"�?��6�V�QB�Ž����[�1��q½[?nɼ���X��<���Ц�h�_㜛Ǒ������4����'a��U@o�(^$��St%G����|H�Ä	4����%�-2܇b�OeVP��p���)�P���ʄ� Z���J��@9zݫ8��́��D��D.�$�%�	����C[�*8�e$�����\�l ���}ʾ=��Z�M�0<W���\rfW��7����@���rr׮�Y��I�/C�x.З�x<$ځr!�.W!w�g0dlei+�P�=;0��jԧ�|e�ٌ�x���5��G�����/���kb�6�0�i��I���{k��7X!_��+I83�e�u45���zݫ�d��&7^doߓ�X r��Y�}!ް��G�Vd�+G.���S��f��G\k���f�����a[�q�`�T~z6��w>`à������t�o��RU_~Πw�+��"D	�\���gY�Cu++�NS��j����Mi�Y��l�g�²N�T{��$G��db#��x�I@�?�b�I����z!q���p ��"&4i�?���&�mρ2��D]��~C6������{����χ<@�2?�Hs��(�Y4����u��4�J�F=�~�8ͤ�Qe�#�5C7w���������P�$ �}���PI�w_J8Gҟ����9��FC�l���2 ��3��)9�(2�c�"`�-9���T���/�x@Y� ��{����)U�q�9��b�b���j&�h7�e�4^3%&��_7���/�O�P��l`����.�Z�����h�H�v~ʰ �[r�􁛄�x���ܿ�5v���T�XP��n�9�n(������D�ɗ^#�ءKx��l�.�el�]¹hJ2�W
�\�L��M��n��A���3h�	�2�:�L}?~�X�{$FJR�,���`�佲P��2~����n������hބT�u�nѤﶼ��u�ihU7�]��+��Տ��'^Mg�h}���Z���tÌE��IN1S0w�/����o@5ւ�W��"C�;���L3�]��h�%���y�m������&��T�y���p,8�Qr��/N��Sƺ�"oj{��N���Dh�!�8i�H�|�j�R��q���$F-���=������l�4+�1�-<&rbi�p:f�uY	An�"c�f�(�b� 8��w�a�z1T�
��ɓ��$�x-2rmt�_Ǡ,*4�
���K�d��\�V�wh W]L�J�F�|/S� �~�:����_r���,������j(?Q��^�8��P6�j�Wi~��mr�GĀ��|��Rv�l(�^�n�+9�Gv!�#_��;|����.4�D{7�1����؋퍬����f3�O�
c�1RlrTX��������:�0�5�n�6��<U���� ��kH(���9W�M˜�Ek9��� �e*z"�B������C�V�'��
��+�g^��G#��H���\��"����,���A����:6�0�dY�g$z���~lq�}�n��D��_�	E��F�����	��RJ��4-�B$�8�A�!���"Ԇ����(2N(�Y~�ҕD(�����^�����%,�s̀y�C�wL֗�Q ړw��A�E0:���(c6{�S)x�g >'C��0�
��%�P\нL̰n��ԉ���vr�T&?�3s
y�MK7(e�l/�ԌD�[�L��AlsgW;n�H՟Kv�UfZ6��)�g�Vv)�ɊmY���?ܵ-�Ti�>ah�� ��(~���\����ދ!},�Rr�ͬ���0l-���/	H����C��uE����Α�����~5!��$9#�],��o����*�kf�;��ɺTg\��h���N����lr�,�f^'�~��_j�k�a-��bH��� `C���܅���?����OC�ʅ���ǱkԫM�_�[�}�������<��B�<��3��@�w�|�����
(XP>M8e���B�\�E�TW}��q˚���]K��S�%mAgR���5����Px�۞���=H�ZsIFOhLx5�ܻ׭�h�O�O��!"l�A58��[E	Ì�#�r沼�֖��<b���X ��5d�4���6,+Y����@��׶>͎��v��?�hk���q&�W��p
�������S�;C�G������
�[QG��\e�M�qoFu�#(K�����Y3�*�G6�����h
�}z�k'����)�_��]׶/���� �;jD.n�B�*q�	sc��FE�#�X�p��8����4ڶ0�����d
=ȀK�^@*��C&����Q�H����$}��.UKPb����6��,�<`q"5�r�J���3�ɴ�
'b�hD����`���v�^����cI��ISWs�Mڏ�%c�"Uu�Z����
����k8�����$���w?�V:����ȴױU�_��*�{a~]]�f%�� ��O?J;DG0�,w���o�_�L���Y$`HU�_���M���v��v�����,_�;r@S��j�}�Q�T>BN�D���O�j�<.���3�ֶ��ʏV�U���qa��	�t���s��@,���c��h�.��F�w�탗�)@����&�}��}�%G^e2�Ӗ��.��.||����`l��_�FM�,|gQ5~�n3�'��T6m����st�?d�!�r���v��n�8 -ⰗU~�^�Ez4�LB�eyE�)S�cO�!`;*�n_�'��������؋�-��U�ߧ��ޜ��!��[H.0��w
��E:�"w5��A5�\A��N��6��O��'��2gy�N� :�N�c�t_�7NGȦ4&68����v��f
��Cw����Q<�􃜘u@��5rr�H�yޱ���M*�h��#UM?���n��TgR��}z�V	�
]7\���vIzT�Ř�u~��ϜJ;ZUH��N���n��6�`̋�EP�\��Bk�k�n,�xC��c�J���Ҡ��+��
�ܚ�N��r��вk�ۥU=��q? #&h9W�}J�I��A%TqJ����4d�; �>?$_��qĔ�,ĎH#�`��l ���C��$��e]<82l�D��X���.P��
'bL�y��殭�� H�#u�,̻�RI�ȷC���*&��#��픷�l�KR6�u�k���ή}O� \��:F��|Uz�(�m�q@+6?��E�ܣZ��h��&+��~����V2����2 bݰⷆS�̤�8�Sm�aN�mHF s���CZ�����4���UF_���T�g��q���clT�#z���xN�[ �vY>d+7D�"yi�#4F�I��3�>lPTO`�����.�2_�N��#{�!�0�Lj�>�Bc��j&#�ԲW�0��.F:�؋�L��JN[�t��9Q�r��5�'�d�Y�}L�%���U��Q�&�Io��Z������,+���vl�(&�؀��S<&�
��)����n�����
,�b�J͞)��H���}e�Us�	mާn��[���$]o�ϣ��9q���W�zHO�ͅ��f�y�ᖼ+��qn�дa��q���!͏d8�b7�����vTC�*�N8��O�Ǭ�뿚R��H���s���Z��i�Y��V_��qon�KOI��#�)�"��qz/�b�~0g6.O����,�0F:�mt���aj��S훾m���>��y���h��zM�����=A���v�r0�g��H�Cv��(v�7�D��B�!N�Ŏ��u$�6� yDr��Xewg��,�j.��}�(,����X�m�����t��IFL�ԁd��TqZ��	
����f���t@e1M�ス�͖�8�[��4k\���V��,�("v���x��T���N):̥�J��*K��oՉq5�S�Ď����T��?���jՒ$�C��Ր�"��έi�M�`��`ai�x�L�d|B�>�y����������z�cj+��N���0ö,/���㝁5?/�O'���r߄l���BR#�����g::ˡ[Q��w���=Z/��d�� P�?ҟ��d��B��!��	!t3ˌ?���y]IZ�/���2��#�K�`�/�mV}e����X�$��|G?Ӗ�o�Vs� ��\IV���PZ�6F����6��!��㫦�bB�\�u`6(r&&��#�rr�*g�l�,�;��tҪ,:۳~�Ȓ�K���%�n�UJFl�1�S��s�3��<�-�_�vw5����;kǙYd�eEHT20Ȯ�~~� @<�|�^���( �B�lnޡ(��9��ȗ������zD�,zX�8�2�zsc�m��>/���S���5�pI�Y�U]�NL86� ��̉�����v�a-M�ٸ���[�62=�)�)X��w���"��[�����D+�H�Lz��N�_ͣ��&sk®ɞ��.xw��p~�bU
�U3n�qp���^21/�y/tv-�e�k@3^t+��Y�	�ه��  ���.���Q�+�-�4bEd�[WI�=��QlP����9��l���V�97����%�����W��O��q}��r����	[��@ ��T�*ف���#�	�N
��ű��F����^���A�g�l��nT�vZ�]�1V����R�H�Ȉ���/�U=v���1ɳ�3G���$XG���KPG�Qd���M�ˋ�қZl [d���q䭬���54U����²iwtb2~1o�/�����H�����_�DΚ��6�G����I�b-;so�=��b��u&�À�<׀�(H�ǝ吼��m�^�[U�����;c�w��l}�\j�(�E�$��КIy`"4���J�᯷�/�z�s�~��(�����j�k�YJ�N�,��-.�Np_��F�T�y���_�:�[s�|w)<����vj&���kGA e�h]�X�%�� ������h�*����݉�fP0�\���M\;s�!��+�����IN����*�$���[��cH#H�X�7*����c���_�M�����UW��Y�zy��!�k�C�L@ye�P�i���U�57?��i�f���k";ɾ��#��}���o�?��am=�NQ�JL��{�EĮ�������9�휓����;3�|�H��W���s0rK��*Yo)����U���0�m��>̫KO����,B��^F$��HOh"�0cN����jyަt^��Q���F��eq�
�K�pa�VΈ�Ҫz��v�Sֲ�	c6=�Jj��3�
�����o=^����h}���J-:��?W�y;�l��l6����h�;��������n��Ѝ7S9�d�=�� �*�l�r��*6$�'��2w�?-����.�$M�����^´	ƫt�-��de��COT����؄1��(���.Q� X9��2�2�gX0��������&/��k�>�p6���:����w��	�B2pjt�Ե�߇*��b��K�V�b�&j&��-�j1�a7+��0N�ѯj�7fFE��%4���͝�b��
~xz������=C��GYFX�>�C3����j�xs���hGMh8�������-R�eQY�@sYǹ��oh�#њӁ�îl& ��p?���\��)�WޓR���3^�m�� �O�i?<����)�� Y`��Q���y�SZ����tne�����>Rvd�~�Ԏ圡��uCr0Q��R�mz���+PC�z:�i=��"�Rؤ�c@�fa���"N�/�_Cc��	��"?S�]j�JFx9X��RaJ�R��Gk�׸Vo�����0��� �ߧ���$�M$��X���I�zz��A�^����H�JN;�?4��c&J����J�>bxjWv���V�5�%#^D�ƻ�l�,ي�'�XZJ�c+�����SkT��.|�i��x����n;��&��9��z��ID=��Un�:3�=#���}���ٍ_Jtg�4oM þ#�b�L��n��;+i�p��HnDhK�G�M뾐<�1O�J`R�jaƔ�����VCm��;�|8W�5��)e���ngT �&�<wShj�q��P���9�(ⱟ��G�0�O���j�,x*x��㐈?��{�/�+�4^��a��� ϒ�^a�};��o�D{��:�PE��� �Yl�Aw�0�y���-��D�)w9P��&�
(�r�ǻ0R�l�D�]�.�+�W�O�W�b��ė@��`r4�,?H4zcCn�r�JT.��`?��>b(ZR�x�`�Ƹ�p�H*<M�i��>~
�2�r�jϥ������:x�_�5���u�����r����!L���P"V����%G�C�IW�1�!3�#���tQʥ�����x��l�d��3o���,+�z��ЛA���S�Qx�!���A�i��71�?U��r�U34�*�!0�c��~me]��%�"��Ӱ�h�&�?Gt�#(�i����E�F.)$o~4�����?Y���p�zS��S��/y�R��e�q��}I���=-	&���& u�]�?���ޔ�t���9I����}X�G�J��Fi�Q�\G�2wy �5�_�*L����{����G1�b��:D�C��j<���CPˋ�s��k��]�F�������a҂����;�0%V~�V{�7r��M��׾g��op�D^7�Z��q~@,h ��+�]`��;���܇^���!��c��3�VE�<1�s{���$��[�2x�*�o����Or����x�m�<��A�(�]������c5��F<�S�B��ss�oh�i��qd}���3�_P9"ؐ�q^�iu��^ҬX�K���0��������v���N�V�4mC!�:k��T�Ne(�<���9d�+��`��j#J"� �D�ݺ���-*����{���0?jšޭ9dO��K����1��|O���7B��h�FK�*=Er
oz��'�2��V}O�0�n0�(��9⹒P}[Q
��ġFkW��9b;:�hf �߱my�^�)�ڂ��i0_Js���
�@1Y9m��H�iEv�wY]���H��$`��0��I}�uSB'�=��]?�"U��{�����W��i�4ES�ܘ��J���<e�~�xv�ϰ�r1E9����'+�W ��"�
+/�p�O'��`���=߇���N�H�/�++H������K-� 4Q�1�%[m�Npښ|����0M<h���/Y\��4Đ�R73J6��q��2��pw6�G<U��j!}�b��5�A�>C�L��L�5&|��Y�hk�;&=�ǃ*4U�4a��gGP6�r�%�������θc�v7�"�a�Ӗ�s��ɱdI@���[�ۉ)�:�.	���\�6��%�L�9a�n���~��l@�>��I�F�v���`��
�z��|.x95Y�M�b�n0�o��
Ru�S��{^�|�fLF&R(�g��o����=r�R4+6��,y`��˸�l*6~��Y�X���s��/�а�)�����H� ۼ�I�6�6vj��������\�Y�I���x�j�:pkH�����l��� ���������2j?J���Vn2.9A���k\�<F�B�a+���B"��!\4E����ػL�r|K�]�Pnf��{���7rh�ω=���?r��]CHȥ@�׷(�3t�E�4b ���*��Gd�D�ꖡk� ��UQC��̭:����Onq0�R��4�GƧ�dM�
U0ض�휴�9⏀lR�4�~�_u�]�m�Z���1[W��|��K� \���=�WN����әV�!�^��̸�:2:J�6��{*�x��{��ͯ��fɋq��a�KK�n.��ÄW?���O���8����1�FR˰�w,��|1W�����i>,C�Q���@IϤqS�����Sg&g���o9�� ����kG�=��,w�ݠ�>�S@)�%�?���F�=�,�I]na|��y&#�@����}�Q?��Wo�H��w�2����{��M���Y��2VR���23�T׽ĭ	H�*ׁ�F��.�S��s��DN20[�MH���=ٴ[���֧�N�Yћ��_�p�q�>;��9U�[��y�.γ�%���Yh�K~�З>lN�z-(��x���_kqOx�ĭ|#j0�k��E	����&�Z��G��Bo֙��kV�J=x���q׷F,Yly��k���/���c�Л�����$�P53)�!<I��r�5ɡ��-W��� �����n{�f�?�R�y��l�c7,%��t��3�ek��FzmJ���EZ��b��g��J�>���q��>��/��a�6S�RՌ�R����D���'��T$
7�bLv�� �4D�2��x��T�~�MW���r��\ʏ�YH�ϝI��}����L��?f\u����C�$����`|r�a�/��P�B�WV��r�m��7��@�oB�0Z|-�;��B��ח͊��J������F�sK�@�yEO��?�*�IR%1%1���[�=�
�j�	?�X��G)r555� ���Ձk���@�ڽ_�JCj�=�7Ƃ�A��6��Ŵ,�]��9�a� 	.��qD"h�b+b#�VoZd�,�����뽋�Z��E�����j#>���/������̾ �VֿN��SR�F4&@��B"��z�;kÙ�=��%�ݶ���A.��F������X�ֵ��5�w���4���F)�<M�@O�g�.�Pc�p��՛�0�D����lkQ�Dt���f���E1�1a!`i׎�����8���h=�8o}�}v�O���"���z�N�r��ȿ�
���s�r����?�y��@[I8�Rq�5�4� �S�w�(o@` ���Mo�@o����Ö�)�Ko�wx�nfb����=��o��l.�Ȩ ����-'E.��7�cwfIG�0/�B�Ja���J(��nq��g��P�/��i�<,�RH ���*�|{Q#V�V��9��Al_�k#��p"���NAkO�:!f�z�ևC�I�v (&�d��h�k��ԝ���y?fqE�g~Ev��v϶�=[�H���ٚ� �@�Y�����#� ����0gd-Z^�r\�64WQ9�­�&����s5���fv�zk�-m�#��%�� �93�8A���m�[��)�Y���wǻ������e�u=m�「���h��p�]��,�њ\�����B1��`�Q���~w�z�G�Vl�'�t �g) �������){i��i���{���_s�HL���Z���A��Jn-e��{h�_��(��6��Ch�E��]��)| �S)��=-�c�d��F�w���j�a>�s.��tG�ZJ 	�*���5��@��sj�?
��?_�����)H���%��L�?���N�&�y�ee���xN�޲�9�3��8�}H�T�eS����
�`y�{cgxd��0��c���
�V,�D�5�k��.��e3 C���>�^���z��̬.4T�hS0�ˑ���
�@�t�G�0f]͍�͗g�G��F ��=��J��Qd���۰q�{?�'N[����E+.qZ���p��]!�^J��W��6��yc���H��]�7)`�cՋ	����E�������I��T��Ȍ�J�1@$�}@�:���F�K�me_u�A�.�]+r��4ET�s� �0���2���2x����m��`eʰ�#��f��)B�fQ������N�A�2l#1J�]�p���y�u�2�䇣�����^/Qk��TW��$�h6H�	K�;��d?bA����H�%�IZV�1py�tZ���_vW�_8�cq;��[S�QE�qiNK����<�)�k>��ᮉ��0C��IB��R�!n�=�%��'�9�@�|G�!�N�ۺw���ܒ�wX���P����$�RB�B�)��;��jX�/�_��S�q���I�.���v�mӑt�e���4�҈R�ka�=(�u��o�8�gfS=����H:�P��y&��j��%�ssd�M�I�������6��B�L}��3~�gK!�!s�ۭ1'#����l��+�����o��۲/�a8^U<؆gů8�6�\׶�章L��o�1����S4�\3�7��m�):��d��eE�j��Pوc-�b��Ũ�/�D��tț(V�������9j���j�s?.{2&M&�Nhx�e
�냇��dI ���HO�� �ݙ���5�H��Eq�ZF,}���"Gegk�pf�͑�K*Ѯ �M|��+�0��~)���{�����U,�Z\�ܭ4�j<|��J(���e�j�M��{�3;b;�l�F���5֕�8��Ġ�q�Z�3�jH#1�R&����p&�}��9���u�>d1�/csݻ�3� @5z����SF���E�޽܉a��ôD�����ٴ�4�kB�ezF�G1֩��(��g�2u��
�nF�9a�aPUϽf�t�;���)���'3B��D�<u{Z�9������=�e����Jn�+L.d�?��)�myԤ�u��gj�Y�)��Y�Wa8G��V��&�b[�������ARb�����8V:�����,xq�r�g$*��#n�� ��Nqm�E����sA�u7�%г�9�k7��Q4���W���X�w�>$�Ԥ�j��l.���T��^�VgGg����wxתĐuߵ��bɥ���d����ɐ-�����,n�i�-�4�m�&�Ps� 1ϻ�Fzc����o�$�LK�g�'=��7 �2P$��YQ��I?�)�����=�������C�[���;08C��|a=54�U�6�s�xD"4-����7�܈�>t��F*R�������R�Ȁ�Z8���m�qZ��8�y`[O'�������Ϭ�.S^Xl�Z�]�B:m$=��C4�T�Z�����l�Te������5�Vb���?����#
�g���s;��ꏗ4
P�C��2n�A�S!~V�Ш�?z�FE#b�t�A�>"7�{�|Y�F�sn�� %�Z?C3�:���\�:���]�B�qQ��T��ޖ��<GӾ�ܾ�*O�F﹩p�J�����C�Q��k��f�}K���0h2�1�������#�����O�s�E����.\�$��@b�.!�f��T�bT����H�l�P�`,F��HW#aj��+��|���{�f�Hm�c_Ӎ
��rSJ��E�,�Ω1���%��o����x��C!�-��C	G�c���s� mL����"��^��&;��n���[,�T8t��x���J��_�V��Z�z^) 栌iBf�Rh�g^u�����{q&�2\h�~(��@�g���K�F8��E�Y����}��To���y�#��d��鮃�'g��~\Fc����?�y��0������Kpw_���POֆ{Y���!���_ct`}�Ѐ� ��l��,o�MP���Tz�?��`=z�/|l�ڴ-w`� �2a�*�� ��H��]�d4�ޣ)����<���Q�a�~����X�ɞs�7I�B��5��S��C
[f��8}:��8��	8ʺ46~m��vD;���)�s��Aᮈ%������x^�q?&R�,&Np���Tೋ�������^:���bK����a\���j�/��k��Z�.�@���n���L��l�.�NvR�\ͤ4�07�>*M�s���$���b��~�a��ђ�v������p7(���͐#���w�<�wo�"�؁��z�J�6����������$���t>堛j���`��qx��������6�G�~&<�|�k�}A��L�5�_�"xʞ�uͶ�����k�vr7o��M��woG����d@���f�{�w8rQ�#_f�HN�c��X�cq�y�?-����/f��=qgW>�X<�8�:&��������8��8��*��9:P.��BA�A�ylN�v���&9���$��Me�5p�ddÜ��R������x+���0wxl}�{1U�"9͂��-����F�{�0 ���/�`�1�e�r��_�6��l�K�'Ϙ����4���Q���3_x؞OiE�m'`��o.|d��R>��H
"��#���(R�"�d��������|<�kZ�X��HN�gE#�i��IPXs����&XI�ձ&�0b<ݤ�Hl�|�Kɨy�&R�/PQ��ʨ)����.�2�(��9짃ͤ�aT	U?��U-c�r�k�ȟ��h�8h��!6t��&58����,)Xھ��7�1�Lf��U�A�r*�����i��g����X��q j�$��j�+K��m�ߓ�dhWmC�jT��5�78��� �m$==��O���:�3י.�V����ԇE�u݊Fp�cǋ�J�<�X��a�[�>�Зr�q��l(Ş��H�����S>�G��V^��d�~�O�.oU(�t�B],ߙP|Z�P}��htt׵�F��^�ۄ�m7�fIqK�*'43��X����ɴ�_�D8��1d�Q� �qL��
����/y�X�K��}���/�7�@l�+����"�Ck-H��S��Ÿ��?�g׿g���Q�=��i�Afv�X��� AZ0b1P�z)[��d�a�W6?�Rr�Y&���u��	os��o�~R�t��f�s)��#��[�u�VxX���S)2�֋T���
/3��S~(Ն��:�|Ն!6���(1�R�鷧myZ�D�Ͷi�
gz�S5��8�?�}r�5F��2�MI)A�:�C�[�<cIak�����$(ݭ*��_��E��K��f�jU{ ͔�;�a�2&mI��e��\L~L�Ҡ���1y�ެN�ED,#�&A�I���cp5W�3�R〇��/+cOD���e~�e黢&� �_����ܔW{�2?�gr0� g�κ�7T�O�},;���X�ڥk���9]п�u�,�L����"r��}��\o/�odԪ�ދ��o;���v��O�g�8;�5�]*�d#�0�@V����������vs�h�8�Ú 3ŷ��7`Z���||Q|�u��
$�֪��w��4�$�nM#q�:�mG�ȅTs8
�p�N'�2[W�q����Ȗe����Ah�xg�[	��Qb�V;8���2��&�E��fI)(���lR���I���<W�H��>�
��D\�����R��
A�7J`݋ٮ�>w�{Ƚ�=�Pw�m�
dV;tG}��}��x�ٙ�B�)t�M|��7�蠧��X�&�O�ǰH�2�Yݟ�{�,�n�ΐ��Hdcˌ������(SU��Ȑd$���0M�0^0+ų��S�3���Djw�M�������5^�#M��Ktf���9��'��S�:T�WD�\#�P{$�wc��m���E����%{���M!��p1�c�}L���L�ʑ�̐���ӵ���g�j��M�NaF[|��8��-x����iPU�"yQ����NJ}�������_j�w���e*���`���>uh��1�2>ƳE���JbX�w9-�#gAl�&�3\�B�3��%v��h9L�e�����N��"�O��z=�p��i!��=*t���� �J�2��)-t��s�u�{��:)��l�MBy#z=��'*�n�'�D
�TI��:6���t�67�ԝ.�
�A�9 Ɍ;��ͼ�����������&]]�2ϗ�r�d�=�2�&X�J��~`��Wcz��oF��g�<�Ŝ(��;�r{ ���a���[���`@U�Հ�ľW��|�iA�m��g���:H����j�43}H9x���{��sl�ӂ�\
1\'ww�� ����ۮ��������Wn�I����o��Q�[�.�!Ċ�i�x�|K��֨{3��Y{i��44q�c��%��W�Oiy ��E޼mV��z�C�������ήB5z��ψ��l�e�jMCg�i,5�M����9D��=\XhV�quހ��&�c�b$�&�`�]�u)��Θ�&@�t�5��k�c���`�"����"� 
�zbiq���P��sб�Ѭ�d�O��¶��]��bu@�j�ՊXF�E�?2���!�,���.\�<`G�!��WA�����8�i"u}���H���|x�r�Agzw��yi�����"��M(+`����t�_��.��U�3�8�A��i(��`T{�RR��۽P���\�����l�.� @�w�ҹ[��7;� ��)�Pf��T�+򸿅���D E0�*�`
H����U�Tn��'�|�П��+}ǕbV�  �Q�!�����gf���8�S��V�1
��U8n���GDd(����\�Ƙ�j�Ѯ��M��^��`�\�Y[Y�:	J/��*Z�U��.H �I�7��X��Ū%�@*�S\
I�<8�4�k��~�{H?T}�~�]��uP��x��26c��7��`Sl�,����~�B�u�}�h$�F�Sɠ�@qo�ⅾ�aQ�H��g *�����:��漻�C!�@\ɱ/��{E$Ro4Bn`,}u�=2DHhD�pu����^��9];�|m>�B$�P�AִH(��윉Q@ 7Z�B�xz5�H�v�����Z�m|R4��uHYJO���JaM��+n�77e+��0D�Z<s�Y]J�s�Ȼ�P�	�Jn"���oy��A�4����P=�Ϣ���Ϡ\��5�q|`b�S5\�G��n�xȜ��ҟڷ����n��n��y ���0dǛ���2�D)��g+L��|&Eq�j3�g���.V�y`�1��yR8�9�]��'�h�ɓ�r��N�� C��Ա�bc�,2k'���U�	 �ٻ��u[��y�j�,T���[����+�� �{������d���O���XY���bzl_�� �����m6��!x��˴�у�5�2���C�Pd�C�R$T��(P	_��U�.;ܱ!N�1`[�쿠C<c��~{�@���":�Љ�ޡʨ���Y<�c}8�S�eZ!�O��<)1�_��n}�[����9���Cک��#p.eeb@�F���,�?md'$��h�g�7�/K��\��,24�c$,T�:x�)=!g=Tn�X�z�T��1�ݣ�hB��x���ζ��K�{U{�*ȳ���V\���;Z@�+�%y�91�spt���c ��c�[T����h�]�a7���P����o�����I^�f�_�,#k ��+a��V�+2")���wX�����=�@Gѐ_u�2co-���XfZy�4�~������=����V����"����z\��jǑ�*G~j�b$k%:r���'K����(_�ݩ�/��A��L\x#( ~��.U\���gT���zf�;�R�ho{^o�D���0����{����@��2��x /U��)�C8��mTA�+�'��������J�3p�\HΎU/]���(�k�e�/rܪe`�2���Pו��s!�]4�Z�Mo\{D|b���>���L2tN3��ڰ1Ϻ��[�d�ڙ/��F�,\��W��W@��<�_�E�D��V�xU9� 2ʝ-t�4��	�L���|}����r�sߑ�+XNO`��_����հPo�[�V��E=�"I,9��c�V��a%#��2���Ap��E���|
Q#,/�1^e-�"YR��j�$a�GnU�F�UU{ʶ�Yc��4-~&���>g�"�(�W��)�4���x�e"-�Mb�ߓ,6T�ʭ�#v;��b-��?&&�;����\�������,@O�u��Ɏ�t��(��K�O)>��*,�M��X�s�)w	x�4UWeO�ē��%�H{���)Ż�̏e c����wr���ȭB�ۋ�x?�>A��*{�+�W���X~��#V'I�~��<Jr,��	6�&e�����}��WJ �H�{�q�9�XH��T���lcq���V�+�Y����a74u�܅=N�W['3���O���\�4'�O�i��{��t�ij�w�e�*�q���Cm+~`J�nm��V�&T�Z�AM8���C�iky�Q��<��玿ˠR�D��L2�%�� ���E���/�:���hѯ�Y���5�n�ג�ӆZ���蟈�
ճ�B�+aO��!��������C ��hD'�T��@H��Y�֩A���3Fw�zo�oB�
�&�^�v���?�.
Y��?u��4}�|J^*At� G�j%am6^2X�2��HqF��j��ҚCp�[�,~� �us:PV�/���X�'�o��Y�B�~q?j�!e������_g�9��f#�
�r��q�s�CGQH1�)�z�T�]ؚl)������]���lܞ�/lWlb��!.�� _tC�G����B;�ԏ�:�Z������"�N%�=?�ǣJ3�"2Ga'J��V���K��>���Q�'����nsL�Raw�V��8�u�3�����b"0c���t�
�%�}D�
E˺Y��뭩!eL刈p3�H���Scyl��(7�3Dej��QJ��I?�P@Vi#MPȌ�e�4���O�����	?�g!�l��{ͷ�4!@+Tqt�y��R��P��b������@¡7ܚi'}�Ѳ����~�6j��z y@dBW�9��088��O������5$�a}MW����>��(���%�0J�B2�6����aJ�GkU�JЍ|q,uP
Y��֊���L��(� X��?��yC)
�����0)3�C����B�[�[��m�����ֲ���(0�u�8&G� ��m�;e�^Y�ڼ�t�1:�J�B�ܷy ș7���,����3!��r�������2��G+�1!p�ܽ" ��-! {x�y\��&�uG9>F�f��m�=ȡ���_eTa����`Y]nc�ʧ�F>�A��l�SG���D��2�ϛb*9�� }B6�Id�g�F )?��0���iMc�jXqn��B��{�ޯ=1.�:�ez(��)+e>�&���O�O^k�{�4Ks�*�CŅy�ڼ8fF.p(l�7����0b%sI����j��2HIi2ߩ���;՞�0,DY���7~u1~)!9X��FT�	$�k�ۜIge�f��3�>�*�;}pZ��%<ӻ[u��x�X�Q"�J*{�D\�׉v���_j�����3�h�GR���NU����2/?#<�I�Y�Z��z�S��Y=�9�n�A?���)r �W�l1זذ�iU3}����DRn���H�AX�7�d$�A�5Ʃ��S��/���Q�1çw��!��=�C�+`�̾�Oi���{x�0�a�I�t��k:X����$��P=I�4C��NP��X�EY�`���cϗ�le*s3]Ufטl0]p�A�����ƹp1���ͅ���EK�}��ѹ�e��g��`�{<DM���~�D���W�m��qA]���ʜ���a�u�20?��a����<4�b�	��X�n��C��� �>iⴖ�A��Y�}��Gl���-�^x8@|-����D	a���z��3��X������F	��#�֨������y����G�{���N�烻Q�>;��#H:T�;��1�u?�!���H��I����~YEv��:]��m(&J�.ɓ9v�]����E��彣~My#�SywK��)1��dŁ^n@�di���/�*߃��SV����A�~k�L#a!+��[�?a�J�զ�W^rGub��.�����=����1�`��"ޅ�T����o�k�"S�͒�w(�9@��V�s��=�X��b��>�e����	,����'�Nc ��F�  � V6��v�}VFM���nЕ������yڇ�����Ϳ
R�q���ɋ��lD���[X�LQvav�����Kq�<-�Q����,'M�D�g�4���5ZņtT��6V�^{4^��7�"�e�����8C���\�s��q��&}7n�4�JKd asEdRO��9o�^Th ��r�8n���fv4p���Y؈���X
�ŗH)݃�� *ݓP��h�w�*���牏~Ư��,d|�s��g��������3	|��"T�߆�x���I �?����+}��t^K�Dam53���=ۍ4?s����׏,�c�G3ޜ^H�}�(����'3A�Ra��:eݖb��Q)�o�{�_�H��{ʭwǩs�m�k�A��&'@m]�zo^��`������[�H�x;����vq��ö���S�0�ԀhB�@Mg�81�{O�u�zpV)ޭ�< �X���C������$Pыϗơ����8x��8�F�e2���'�N��+Y8�rT%k�^��^臠ز����	���m>fޫX���꒘~C�@�w&P1������o��Z�Ki�8�Ƽ;���๋�T�!i
�1��x�l�$s��x��ǵTޕ=fHV��մ���<��HN��X��|P�~l��-�<>��xn8%+�{#v�kX������@�.�=n�_?#\����;8Vt �賤늊��<���\
{4׫�G�g�@R�a$���`�8�|����AAX��d͒�H����0�f���N(���UF�{��[�Q�Z�Y�	�:���lV�S�+w�x��3�,��liu!�"��o�݇�۫>�%tﰛ�C=�U���7�5��A���O�ҧ�%�{��:�׻O.�,�*f���{�R_gH�ԅ*]N���V�',a���V	J��T�:��漑o°�2t�u`Ӗ��*W! `	!�]�Թ~�?
M(`&;��/ �IG�.�!i���k�n�e���?�S��8@�'�y��"_�]Y�E�= L�IA�x�_P+0�1��J�9���cZ�d-NѾs�e�Zd�j�q������)�D��P���Q����p�%]���?*r���-
��5��A�Q�j3Xp|W�wr��އ�����z�}�P��H4Z���~�N�W�{r�)ě���_qg�5��V���]��ls7O�b n�ྖݽ:#`x�$�i�;���J�h{��"7O�V����#eʑ���.n��2s%�Lc������(C
4����Y#W�6#�NjX0�9}�݀s/j��?:p���e���R�4�,���l�b�9�ڶSs�LЃ8�)d.�_J�e����g2Q�.PG��k�> �Y����l�{=��v�\|�T�XNN]�0����KTcA3�Pv�˃;�4����Z_���,����\zT������.��წ�}�&�+dL9��+����ܥk��i|��Z��KcQ.Y��,Jp36f9."��QӞ��ufʂ�{|�&/�I�]�.� A83a�����F�K�޻~7P���w'�j~Qt/��Dz���i��l��ώ�z���>�.{��۠)�c�R�Z�ݺ��4�mِ�MNV�th��������ܩ��ܶ�0|�e�,�7E{�b� nW��6V<��B#D.��/@��)D�X�sb�$��R�����f��d�80c��j	������{���hu�6R�W�x}(�y��8�*�#{��"�����P�[�� ��|D؍�w���%|BI���߮�f*؜������f<fm�V��` Zy�����V�wZ�L����Q޺�{�H�>�̼9��u�j�s�����,`.�����f�q�`��tK�.�-�S\ؽ6����w/
'J�ܳO�L�z�Z�UML����j�B4���� 6eQMk,Ha]�zŜ���1P?��;���vHc�ϓy��&�픻Sttp�H�lԼ��d��b߉��1$������v�k�wzYO�E5SS���R(BWx�h�-FL���]~�:����i�<�&��?�`eV����FaOZj��C�{���m.ΰ���ݚ0tp\����^aG�5U��4��I̗��i�����0>H�F�?P;3�6�r�X��#�������G����V���t�g��-cU��D��؜*)�B=��x+�G�%='Tԕ�/�a7�Q^pn){G,���=Jߩ�	n�\�"���͕�%Q~��L�q>�'J��X"�.��1O$$A�KP�d�H�٧`���R���5� �K���#���Co��0'^i7��@�X�h�"X�;��S�s�H��J��ԍ�$))����}8Km�[h��	
��%ڐ��"b��缦3���V�"]�]-��)�F%s"��zw����ʥ��`����c�h ��p���������˕A�N>w���#qC�<�.�qar��l{{�,9���-��ҟ�My�ҮW��5)Е�'i��lF2#�G wr?	��|!R�U�@�y~0`<�?�a���6c}����i�P���/n�)d��c�˫(:���m��}�ݲQ
�)�W�ͩ��r�'��#�)6�\�/��Hd�l-�m�{ed{W����$ٻ�^�h>%f�H~!�О1WW=�Ĕ�v�YR}�ث�B�[4������4`��<�`~�ɪ/��)�ڧN��pn�Z�p��)�9`�Nf��N�֗sc7�8���y����̥���L�)'@�.�!�'UH�w ^���|�7� P�̵p�p�Q����Z���T�2�e�{H����A�^�v��yCL�~"���s�WN�v���(և�=غ�0�m�t͠�^��]� _R�l���һ�Tˬ�=X��S�.�S�ucA0Օ��gw������C���;Ȯ��a���ڭY+�s�%�v*�*���~J ^:�����M�eX̷&JtY3��7� =B�����a��W��a�}���=����F֕���P�.p��$�+�,.ru���nrs�(/��b���vAn�"?��{�"��ʷ@3w47%�X����h���=l������H�/��7�k4a��\�WG.�*ȷϱ�Ԯ�-����,��"2
+��$*�K��L�<��E����~1]{��{�XA��T�e��˻Uq��B�Xl�3h٧��~�ݳࡴɻ����"�:3,�a��?FJ�1�x[1H��J�i��` �ҏ��D;P��/�d1��]���6�@��\����"`�� >a�ɮU�G� �:�8�Q�%����������[
�S9�z���:{r�m����&S*=���:VH���C��ۀ�-�z<t�B�:��T���*�Sn��vv"4�A��C3���֦ܲ'�(�t�e�W�?ܜ�v9��Ǐ,;fk���(�B��\�����i�̆�u������g�j�}^���o�Lg�3�>�K
�nw#W�ʒ�� ��V�}�q�KBΐ�"k����:��ͧ�G���S^��Z�'�+0����%V1x4*�z9��`GY���i�5xYu�!�ŁQ����=���0$��,�b}�9�Ź`�f4~+A+�5��!��J���K�n�}��M��q��W�`�ޢ������@�N0�� tț�Qz�x��U��2˗���m��|�+�JT�l�����jZX��/�M5�`Y��E�K$�={5	Oj�����m��_L$�9�i&!�4!_[��	8���2;�����{v��~�b�w�!���d(D槞q�p�l;YO��N�u�����owҒuȔB��}n��*��ԅG�V,��*,c����#�&]M�;�
�(Dx5r
u��7�����6��&́n��r�K����!�m* r=ѳ�z���rw�$K~��f��e���^q�20����^����R���4�
��!�R�
'G�0�+ȌV���O?6z����׃���BEN�r�\��.u���͒^��聐��J�b�)� jZ�@T�E�WfR���bq��v��,CJ�BIv��|��ɾ<fۆ`4��҂�����xJ2G>y��y�>����vD���}�-�y�6�D���2z�O��|�["�����1b_#s�S	$����$$�SS
 1���D��G�Zk��S��\�r��;�.5ZIE�'PB:��؋Rs����o�d� ����/��3xuj���gG��\$�I�>w4F�Ma�~@�xZ�҂e�̔}Nζ�|3���c>��n>�2'�Z2MsL�����v�:�U���]�d8����H�G��!<.��;3CʪqF���S|U��g�F��u�|����^nӢ�C����; ���
��FYK�Ay<�V�C�=9a��pi�O|�*��4�4�:�NK�s��m]b���$\�T�=�~�������+���Q�[���ڇ�62h�h��R���}�:��_�5K��tA��{�HԦ�:����o|!�e<�V�5h�&�U${UT��r8>~/Op���f��
����"�L���)��rO�*K���n/0��4|�>\͆�b��Ӹ��|W9p&�K9���G�C�W5W�݊.�;���	J�ږ8��\�P�$��y�xFO�B�:�v`� ��Z5��ɴ���2�7��B��	��|+7�"�˦�s���ɰ~�Lۭb��b>Pԑ�4�z6����o�*4�S������0�63��z�t|�;�� ��j��G�h H�������<N\|�*����Xt���ccH}�Ja4�s����	1:�lK�kP͙�i�����7f�p����Oe��|v݋�T	�,c��pI:��e��; P���dI�t�:xy��&��nC�V>��C�~�!0��v\�>���B%����Z7��ڸY��T���9@�/����-XОN��/����CV�Ԏrf%�r��-�Oү���Y���P[pC�]"AB�<;�)��<$��g�i�9��=�H�[c:�d)[scO;LU�������r�8��ʹ����µ���ߓ(�T�i�p��5��q I��<D�t�H�<��q�׌�|fw�^��u�(��<�p:�O�}�B��:�*�"�V	�s���:q����܊��NR����Zb�P���SiW�:H�Isfk�A�c����yYJ����$7g�2Ow�¥Tg<�=����]��G����q\�!���Pa��q��cQ٭�f�]H�X"[b(60#��]=���{�T��$�N���7�M��+�_�{���z�S{U*3�}1�T/~�|�&6�������G
��'���*�W$#�ڴxt֩��е�4�?��*b������P3�6�۰P�r�v�	�a�J(��I���nm_�]3�j{_2%S)�ls�K2���}�(s����j_�@eLW7�j� B&�]+<��]H�r#��|Q���Y�	�
�6'�W��,�AA�u�M�|�z����I�.G�k.�������K}��������tk;P�R��O�E���.���ŗ��
%k~�8��4����%�ӡf[J���5> ��$�|�+��i��R���|���U"�W���	I&1�c�Is+ӥ����5ᇐC\�g�"��ع`5743���i�t�\�A�Ǽ���b���]k�z�)=)���l6xP%�.�m�:��A��������^۰�M;���m��1&Y�}uJa\)&v�����5녧�=k��i�p3���*�o��9�
$i����PU��j|PX���q�'Ahs�w��ؾ��z��L�8�p,4e8�k�K��aj����O���?��$K�X�і>^fA�1��>ۖj�('D��"�4�o�a���)[5��~{FE��=��Z�YH��網2��LS-���0�i�f��z܁G7I�i��� �i(x���~����g��앃"_�A9:&�T�������(�%3�k��3�����w�4�au+���H��p#�@)�ע�(�Y�����%��:?6�819~~O�>�a�O�Ϛa�n�8�C��`1�;�E�d@��!j�T["N9�^k	q4nyK��e�i�3�X��O?w"�cv� �x�]��������I��[�e�a�(��UU�B��:�}6ٚ>)�}��uƷ�P &1�֘�ڍr��z�!FJ�=��ߩ�,_�K���/���|A��*�z��myW�?\�V��\�lf�|ݤ}&�p��o�4����|�|>������)�
��~����ɔ�
}ۿLs�H7�P���;�sHT.}��?\��)�!�o2�ݓOQi�u3P��/��BV����uϩ>֎�+9Gw'���k�������VQQ��˭|2�h�^��b��a�����U���Ç�Uwp����������x
a�M���c�8w2��!jm��5�U��e&�7�\Q3Gi������-ɀ_Ic��	)�+`����ȱQ�ˠ�a�Deƈ�7��1�
���	���](�*�e�` 0}M�ʹ���L����i�Q8�x�p�?�tr���՞&-�
7� q�#�u�(`>'?[b����6���a�^x���]O�+@�:�S�.9s��B�Zau�/
��S�Gb}T@:�
�9��^rf���A�&i�+=�D"�<��+ф+�D�A�ƨ��E|���mC1���i���Id�\#dXR��#tKQN
�_�|	��Q�&XT��cw��=`� w�'"��6�YK/R�7���-a|����r�n�;.ݔ%�^5ێ	�o�hB">�?�`w$dZ�lï��t<`��#��}��a�;>-��&�3� �ǿ����󔱦Sx��$v��hk�����s͆o��]96��*�W�A��<�{P��L<��M[�N���rr'�L˾>�jO!0s����	��"�~+g3���@ L1y�/o�5�����@���/� ^�-_z�['����7Re���'�ϧe�5ZELݥ,�D����<��\��,�O*/�'tҢ�j������$�x��q4
 � ���Ϫ�6	��� &i�#6'oZfnn �~�c���0u�
:EsC=��t�bb�x (���#�L_���	psM��п
�9��g��ب��7T9�p��ْ���_ᘏ�/�C�d�=�)E�����\�~�[�c�gݜXV���Ɏ�2����*A���s��P��QU�OH~��k��BWG��r��������fg�=�%e��lR�b�f�G�x͜��G�LPxo��<�ε1h�ϼ08g1n���t�z)�V!lcy�ޮ��=Ro<Bٽ��]��!o&��;!dj�2ϕ,������{����a6�[tuq�+���J���c�as�U�S����A�Z
�P��@�r�ə/Ɵ?�0�'�u!`�˸&�Q�5�ӄ't1�����]4����_�0�x?X�<����#)TF�V�+�.��K��[��Śm�'_�z�t�`��#�͘J�H�fZ�M�L���%g�(�f�dk�&�u�N7
����)����gx�O���58ȟ�� '���I��R!�ڋ�i��le����v�t�Y�hx�j�Zʈ��G����dn*��R�t����=р[�S�)~+��e�?��0~}�ӽ��,[��F�@����R M�Po��rf���?�\��l<���;G� ����]	�HMk���1>|�G�\Q�THL�j���䯶{�Ts�N;RXYV=���![s�LHSӴ�R�x�-��V�a�J����k~�ԗ��U�~��҈IPR\#h�����q�6�bC���M�U�9�5z�t5���/�%�'��Fy%)�IfDmз{��З���P��>�I&*:l���qn�h~Ǚ��}�A��E�P�E���˕�"]x�����5g�k4�4��G��Ne����w�*5:�0\��K�����;�<l�2�Us	����W����ڋ��k�a����Hk�K�0��s�P����nBa>���VK�������+#q�Ҳ˰��DK0�a�!���1�@_o��e�ka�ʥc�K�%��@
t��5Uku���� �a�����?��KZ���g鱃�y,���e2�G�X����2��_s0��@��LE�ٯQO�T��!?ϖSE�n�6kR�4��]���"mM+?�))/ ^0]���@pm-�z2�������Ж)�Y��Zh�ڵ��5Tr6�y�r~�Yd� SdUf���v�F�]�lY�'W�u��cY��m�&t�w�D.��݄�5о��*]�� .<�enlP5Ypq�~�	W�6k�D\��P3K��BX���|&��?1y��l�gF��J��T���%^��hef����ݺ=�ة�H�]���ebW���0��[w�V�W�b&��Z���\|d7XL�P��r:��rW!%�YB���g�.f��~od*߷�4(��=/����4y�Y] tr623Ԓt���.ߓp����uY� 	7W��7�m�)ͺ�yi�6SSW�֒��əq:l��3�(��eu�5�-a�M���V�a>b{��2g|)����"#J�Y�w���Ӭ���j���`����G=Q��$B3g�����;$�ʪ����^E�rMU�LF��e�2҄��ƕ۰���Ҫ0�)��={)9�;�5# $���H
ڰBm��ʤG6�(��C��B�(�3�WEe@&K�� ����-7C4f�b��SCWM�]7�T����s	Ui>}�L%F�:�i�\ά���:ɟ��|��7�I��r���NX_0�nԑ���kO�ǣ�kb�NPV��o�hy*7�>�$���4��D)Ф`5| !3c]����-�
Y�C��D_��,�
O�ު0��f��#QM�h�:ipzN�_�m�vh_�����y7J���f)��oVP3@����|!��bd�����
�=�>�J=�x��H
��s��{�<sߎ���,uhl�n'$�z5�a=�<����֞P���T�S�m��F	�X�F;"��y^N�ag�i$T�]ŕ��&�|����(-E'{p�(_���)����,�t�\L|�Į��d�s\jr�l����dZ<�������6����2z�e���+�X���pQ���������7M�3L����W�t���#�o<c	�}�%�I�Y����yZ�?��*n���I����k
�`��PFb0M3i�*���?W3�pn�r�Bj$�ؼ�^�+�J`�T���&�~���2�2��ݸQ�k��%��&����9����W��|̵�'����u��j�̲@N+�B{�Dĝ���>-��Jd�I�ɑz[X$��'��/�1���.u�Z�����]��īY>���o���ks���x*J���$k~����n���xC߾:��.6_iR��� =���\5�\ݎR%�4�c��c��l>�l���"{�d����7���-��|*��0q����ն���z]ʷk{��@��44�m	����+9m2g�C�Q�?��"f���2������ c>��|�f�OU�욯ӑ�m�]��*G���.�xKL*B}�|!��	���͍�{��y?��ڨp�ϖY�#�;�����6v��_(�K���s#O8�%�63x@�_s��\��b�]�0(�l�Q���;n���Y�T��*zid�ƬMc����6�$�����W���?��R"��j�b�f�S�ZI��������|8^�P�hX���u2V��q*�.�o�a%=m �7v��YkB���8�&��%��KI�$~�=�-��������|�������Kt-�H⡆'3q��'�$���6fx�{ A����BO�+��9VҞirez�(z��<ݒ>��&�6��f.�����#xY?�*.��CD�h���U�k�7T�b+�	��vLJ��3�k�p�xq�ϝ���L���J�|�A��G��&�q|�0�$%0T�	�����C��٫����V縤F'��X(��f�0�_u.��1~�%�6�^g���H�S��斱Zަ�I�Q�iTï�Xio�@E�OTͷOz�>#��'AB> dV���ϗ(g�ȞG�Ẁ�KS&�[tT�4x<Y�e��{�05�v@����>�G\���vSI_�1�&� /Ս|��P1�Ҍc
H&)`����?����0/1���t�/=�ļ�N2�T&�]kL���7����x���o��I	��a���5��>�T�$ݿb�0�BQH��Ŗ����'sЫ[�6��薭	�B�������� ��\��|�`�	�;=���D�4
L$ymԒ�c��^�DS��{�5�к��i���a�m�/��2�x*��Ju�|)�]���%VI�X4� ~vH_4���Ŏ�{���r_!�K����#Ax��il3�Q�<���T�!����A8y��ۿ��bZ���	��6w��D��a�z�J�]�3k����^0f�ܘ�~���a�wcmj�(��0ҩbޭ�oW'��BS{���A�D�4.��iL��S|�ȯ��J({?���>����iϕ��9�2����|��Qey�D-^y�!Ԇ��σ��[h����|���-P�3�s������<�������@$�ƨ��&����gx�8,�o�n�\��6��%�Օ>���h�cئs�ΐ �*��=�Q�~;����5�����z�or}��K���З��a*�����U� 8[h�!Sm�|�$�
N�v�U:��u����jpv�y��ܠ!~�3 ����F����ݙ���:�FK�����QMjY��R�I�n�uZb.��Lˑ<D���:��h�$�4������A"p��8��(=ĥ N�s��y,�Mh v���}����}��a1o��~���H�z0��2�]f��5R|���wg��헐��0(O�N%�����2<���M��`�%7<�ӷ��L�&�慓��sH�pЏ�܇��y��78f�3���\(fKBg�xR0�z��}�Bo���c_�'�^�~~I8�4?[ٚF�u�g����𒵂��<�'���FCq�8���Xmnȍk��:�r�ae��_���h�,)�-�����8v�C/�������"hw�]a����N>����H-ա�RV��N,�JZ���E�qP���z����i¾ ��Jo����+����II��x`\�W:5��������W�փ�N<��us{ pB�:��3ҷ��S��R��bD���4b̜�b8](`�pM6w����as��Xxgƺ�މ�	Q6iŸŇ����5G�H�Z�`}P���3��T��rb��C|���Dt� �����digz���P��V��7ǎ3��J
f�-(i% ���Ѷ�<|L��q,�zJ��4�L�q�����z��RUO�7�Ɯ����`KL��������d����wbV|%��P5����ێ�ѹ���~�G�4��_�
���ЅjO�	e�z��H��ެ/eU�ޗ�}���?�e�m�E<s�3�F��(�������� �P��pڅ@ꆕU�C1�O��*	y����������
�~F���@�ʖ^�<��_C;�^���6�1�G��4s�����Nk�����$5�O$�s��2�[�J_�şb����Qh�;T��� -���
�)����F�>
Ք'���f�]��㸑�����R��}�s��~�g���k}�V�1�"�(�eZ�6ϱ�N_�8��x�h-i����&Ѳ��>�| ���� >ޟ�l3ufYY�5��m�!U�7�ߔ�1$�������
T��:d�ŏ�A�?����:�g2��69Q����R��wn�p�7#�K�:iP�p��s7��LF���_)<�uJN�M��Mؘ>[���G`�Bl��Y����6���֛6�D
�ա��_�W��A�S��_�U��=8�f�#�ky��F-�D:��zy����@q(�����;0z�ʯ�ן@��ڳ\�G���ܫ�W:7�O7y�p���8�x�dӯ�I=~R[�R����1�]�+�K�B��.q��
"����{��>�̍����T��|�u�@��6x� %����Yt.��D?>��/MiAS�P�fox�����a)���|���`���8n���.����-K�?R�j'ܑ��dk6K�q�[5�U���/s���晊u2$DPqWjHh��	�̫����olP6ie�"��`��I���c^�|r��<�<�[Y�=��¯i���8�P������/M��D҄Q+�=q�����:q�S.����`1j��1%�Iu)�H����.ڪ5�?���A"�Cs��ྺ��� ���7w�����@��	
�>t� �^�ܪb�����2�Q�����Pz�bs��{�\���W��y����"��ɒ�?_>u8�K;֓ƽ��IoPe԰�{�]��$y���1��/ xl].���n�S������k�#h�ly�s��0�\��.��?#��w<x�.�GZ��DA�(Z�pq���$d��������k�
�e3��Ѩ�f��G�CNy�o�G��`^�f�^�,����:M"���#����E���$�JH��h-�-Kٵ`łT�`)s�y��mIbZRi���|�"��:�V�x�Q*{Q�ҳ3�;�i���	 e��<n,��;�yQ�S5��|H�x9�b�!u����_=��|�� ['���2�N�x��0U\��y1��^�g~{,�����^�pd�z4�i���� ������e�~K�;��R�p<u���E�S�u�%qD�4����Y����Vp�/��p9j`�|P�ɻ���9G�D�b�K.���	��> ��B���x8��7��t�~?q����qel�7o8h��8�V����;DY��
;���}H��C�<��������oe"H����ǇUw**��$Mطu;�8O+��и�IhZ����#��gB�LƘ��X�f����J~�_룾r=v��o�������T��`�������T�Wg2.�]�i��.��	ŘdS"�)�`7�n8ڏ�_~��UU1�Y0H$�n%�9�`�1ߋ4��-J߄wS��#�hE�*k�w��y�	uU!g��p���	�l�3�$/��hb��Y�'�k _6�!�ʡ���:Dn�[����33/VA�k4EP�ɮ;�K���
U�K}&����\�vw��Tm���x�I���T�N 1]�����k�P�8��sX4�M�B�(����ah�]I% �[|����uH���l�OU��M�J�,�Qs�ܔ ��!q���*��yw���k�xM�-(9-���� q��N�"�$��sJ���*�ZzyK��*}�ڦ��o��0g�����@%�w�-{+gQh+�������M����$�'-�4�\S"�7�ܾ+������ͪ�D,�;���ւ�l�����4С�F�%�� ��Bh��&^?�t��~�Xx{u�q{"�>Vo��i��G� ��b��f��\���m�@��
:K�~XZ��Ù$�QcX��V*D7�]���U]��D޿`)��l��C��c�M	�$��o|c���}䫃�����?���ֶ��8�6 ���mZ�n�\0:�p��Ebb���6����<��킏]w�]�9P.g"�$��"���I��X������U�׋㸠E�O����+�TP?$ �<�^`���#�3qo�;V��5� �^���\�����+RX		U�y���h��Cy˒�D��A��Ca�kt�^k�(�����|h�1V{�P�E�+zl*�(�C>�ŲMRɻ�^1�1ǃ��I=��q<���p�Çj�j�%�����#�lmq�-x����;RYY]���ۤ�g���d�} ���?���������^��/��¸���I�G�˧���I���r:5��C��ao�Jd&z=��n~�g�<�f����W �� ��	�������9G<
�`�f쬀��m%}��f��dlD�=���:�[,��N��ZW�gu�!.�g�x�W=ro���@҃�G�����R�LB�_��/x����>0�H)��I$EC��BY���#	AiE��`,�G1������|w��Á�QTx.��r�x}���(��n3�%%<�!�V���3���$�˦�%��7�޵��x�`:S�B9D�N:�lB��a�Ly��6���Λ�+V�F ����}�y75�7:	�l�{�+l��#\���x�e9�~P���
G�"�/�[_<=v�d�~��P[yD�e��yR�;��F�q&�������>ހt�Y"�7~�Z{��"���CFSyΠ�|�O�PE�(m���%7O���kΝե�� K7��[@��7��x	$Ʌ�fi��m n~��@z���ޞ�s�x[-O�,�BF����L�k!��j����gS��,!5M%�����A�NϘ����v���S��5�r�S�{4'��D�
m^29f(�U�1���4Q���y�	4�w?2ؙnI*=�LA@%[�:���>��0;�`���^\1�g{�K^*IB�o���L��N�*Q&�l�?r�ʃ�+�E�����Y81��	eq�s{?Mt}N���0�v�,�n����WW�"r��-�M�nb��|�7��ao?��(��]�O)��8�>Wu�GQ�k.���	�����c m�B�قd�Ui�{�?�Bn����L�������_�!��ff��a�h�^$=](~G*ڊ�lE9%���/�Py���K�P�c���5H-EYR�=����
m*S�F���{/M������&�h#&�GU鉧ִ�
�����6+��l��~r�_EC[�F��>��;��%x\��5nʃ��w
�c�mJ���N
�6��ֳI����S����3���)��|^������MHgՖ	�^ٔ�/R� ���E*�h�uF�=X�N�A��'�Q��+;�Q�NҐ��JU�t�Yձ�r���|j�4����+6ҿ0�o����� a��k�������#T�]gF�/�C:�iTDV3�7O��������!�X���cy�l�J@�tX��v�Jݴ�!f2�&Q��@ @Z.��m�.�q���u{s�8�,�P�Qe���]�Iq��{mN�5��6��׻���-���0��v�����3��;���4�L؎#s�>HǇ~$��㸾�0�ñ�Tu��Z~?tӗr/�M��l<�g �ܗ�%J���CˢyG��ǝ����w<�6�>n�t��#�s�(d-$�.�ff��h�[��I��d�8�Cxpq��,��RB�U����\����S��a�s�%9����gׂ������k/�b�ہ�!7Fj>@j�1�8p����拋����$Ě��p����c<�1�(�?�� �x`ǒ�Xw
�a`��/`�|~���l�+�Z����o18V��$8�gy�e��4�l�z����ihke�WJ�&V�O�N}6����M�<��D{�M�����)�:�ܙ�O�B�q��hH�����|��
����ClR�fΊ�
&A{�9�8���eo̊�9��ОEy%O��cyZa�(�Z�L�XtZd�Ǝ���̦ ��� �p�'�.����Gt~����C���=V�lׅOw� �8Zٙ��lj�P���k�3:7�eج�Q��b�c�(�EiU6B�﷣��.��p���=�*pI��!^x� -�trا�����Q=�ee��N�-y�%���Ȳ_���/�O~�¿�5�r��⍾�ԴQ���L��K'��p�ԑ�=���4*���w���7�c��lm]��T�YDB�+V�3�V{vXRh�a�e�Xmv���@5E��4�)�4�sBK����0,3��s0�ı;B�(�B�����(3��-eӈסp;. �b��eQ��i��I�<5�i�Z������,~�o�ϐ�&����� @m�V��=�~$¾��q����h�D�\[��U.]� A4o�������%��F�)��~D���Yy�n� !q��t �
�F�;	C���2wf�4��E9
��[�q�w*�� ��hi�Y'��Q�?�5���ۈ�`
��4��;���C���e���lCc2�#�u����NI"1��	;�@5=�5���H�s��Jp�F�f���'SPu���.��h1��皟L�P�c�#\:˓@��� �v,KЗtŤ~�ex%T���g&�=��@��H��ɖ��N�c�0z��K���bMe�5°��}E^��*��ش�v��pe�j,����H�I��5S�<����p��ς>ɤ�ܳ{�{l���f��y8�k`��
�I>�� ���9�)W�(r�l��-�%�T���0��y�*�8�з����nY����5�l2%�.�`fMoK�_���s v�>���8ly����Xn_��w?Q��ʁG2������$�\|�alMȉ�k?jwa�%��S��~׽:Tn�Ɲ:�K(8���( -(��b��E�;�y"����)�����m�vV\9����MZ|����-��j��A�#(��,B���,��	��XѸ_-�<Er�|�������<�� bLH�=���!���hB��,�q_�%2(c��c��p��D]��z��:�7�K\���\��?�ϒSq��\a���O�Z������q�G��֏����pq�k#:[�p÷`�n"��o��QY�ӭ��{8H�ǘ��x��$�gU��q�Gb��=}�ˁ�׎J�\-G���|�6��1r-ٜ0�DVL���t��i? ��".H���� V����s7a �%�HE�:�xq��vF�mLx�G��Q�P&�I��>kL�?��r�V�8驨M��7!�L4�V-�����N�ۖ���T�!f\N������\��x����Ҭ����w	�ȡ���(uV�x,Aر`��`� �<eB9K�W�{���f�J��3Y�1����E�_��\ �,��sm�÷�˜]� ���C�\��\�>Rʶ:l굯�=�����nPu�?f7�3�
q!Jk�F�Zl_d3̫��}�� �V�0��ɘ��M1�v�ZL�T\ŬYG�-����U-�'���k�bJp�bO�����(�;_��x��B&o�wX���^�h����7l4Q��!�:4���Mg�0��>��i���@><��=:)�M]���ؽ,��z�y��q"fF4����v����V ��{��$�Q�;-�c�4���j�Q���1~x��i�*�Z����WY������*B"��/ȾG��e��ů
��M���|���.f�<�#��9M��W և�δ$�W*S�r��םjPa{�t�}}CN$X�ط�������w'
�z��_m`����^
DТΤQuΥD�j��K_������s������k�B��ү
�6��zԢ?���Ù>����ha��i/o]s��K�;&� ���M���q�b�i��liC_�?�;�$�C�������5mb�g�Ys��`z�NhMhǦ7k���p/��7#����e���`�d�z�+|t~&{����^�au�GÃM$-_x����v�3�VQ��{�[�cJ�TLi�𡸗ˋ�]���~�΀D�¡���)��Jpm0�o�7����G�1��}�ٗvU*��MN���i`�'����2�¢n`]������z�(�����w;�I���_�㧜uO6��v}�/ @_�����H<��cE 
a�$#��RLQ����g#6����ފ��~\ RRF#Y6�r~�� `:��U�?�V����x�OoF��-��'v��'����Jlp�����=��ޔ��T�p��P�o��j)��l���R�4�'[0�-H��\VP��{m$^��(�'��%L����4�pu�մ_}��cf�l"��%ka�W��)	be!�zN��xokJ�	�7Ȅ{ٕ�b(:�m�~w��iɼ���e��R����*	:W�];�����ݯ_{�����=ϯ/���n�i�eü����a&;�i�pӷ�=��*r��|N���"�N�DK���M�V+0����1���K4W�_
	h�.����/��vQ�}x�Ěz�����<E�aУ��fGB �
w:��0��t�4��X���db�^��Nw��-��7ҁC���$�V���q�u�ī�-����.@�����%%�^Q%2�6c�9˚ ^�������n��b�)������%4�I$#���,!�F��u��6��hЃ��CH��!!�Md7��!ƍ�6U��}���a#���M�wye�����v,����I�C�(�9x���,0�n�DԷV��(>�NR��gwPa��um����vj�M��f.1%�%��g�Y8�4�X���JM>wn��];�����#Ҕ%�Z�4���H�d�e-��p�ӻ��,u��Y��`��odX�#A4��J*=�A �����T�-)!)+P�0����\;��O50TY_����8���� �}�eu�<閵 ��"
����D)qH�3oli[R�9�a.L.;�ғ��H�u��E-P�����+<�X7�S8Ozm=�KO址Z&fLmr[��3�������9�-}�����L���*:�1-���.a�
�d.]�Q3S2AϞ�4�Q��j����7ǆ	�<�\���5y�Py����9e�q)��I��
t�4���-t�	��KQzA	� ��甚������Psӊ*F��H"��աxd��>;���!.���R�`,%^�C�2����t�N��S+Ϯ�tk��z�$�p������	����J-�n�A_���ɽYU���ӄ<�D>- ���L��s��)�ks���� Oܻz���,c��u��*xBwh�ȫ�(]���r��iK������un �ث7�({�2��>����8"ȭ�>������WLsvb�I��j���7�R3�k�=�9+�n��$��S�!şez��!K�CO��i����Q���OrKf�FWI�t��35V�T��x�H�5�],ivADW�εH���y��P��|0�W|�S?ƺcE+KTJ�m�c�;_���%������:��U�N���k?����B��T�˟B��Թ�JY"����9���KۑV@^D1��&�}s��:�V�"�����;0ֺqn�P�o4��
o��g��N3��P��I�(�'�c�S��"�q/V�;#�\(��gg��Ì��I]U��+��a�)lDw�/m��2�g��ϱ��{�b���J�ߏ�puu�g��N	VT�n��4����`�.�a������ĳ�~ˮ�����#�$���ƽy����W�7�tJ����7�Ƈ�@Y���O�s�W�򺽪�/��@���MK���3�e��ΒQ�z��x����\�'զ��u	��`����#�|��T���]�u0|�m1|�S�<�A�C�
|��6̤S��a&�"t��WIK�
3�Lp���>cB�+`m�}"z( ��8H���y2KS���E�"��ne.�b���O �ȱ	S���v(\h0�o�ET�n�3���8��/,�>t�~�7u,�sT��`l!���"�8ÁO����Ʌ����Զ�~PZ�N�#Y�I��z�>	�9=���Du)�W��I��#�+����z#�obT�
@b5A>��~�Z��s詘� ��תH��CN�]��mcB��lɆ��&	�u���|��"��$�rP���������?����ll@e�m7З5��m`h�J݇A������^���G����pI5$�$8�A��iW%x�l���'J� jq���3��)!�2[M@'�]�� (ô�K���&G�ף_d��Y���B�@���!y����+?�"�ǻd
������F��,����3����Z�ǰ��5���;�ǭOʵn��՝�[� ��w��h���Z�t�n��b$�D~A�N�	=u��"�BY%Sk+�w伎` Ւ*��.0�B�u0��S�{�V����i�L�f�b�~
����qBW�@�N����"+"����'5%�R���