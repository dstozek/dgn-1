��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t����j�X�8�����$4L�������}g7l�� *��I������,0�z8O� ��t'�O��!y}_���C���cC&��BB�m����_�2rI~�K0�HR3=�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HCZ�C�Ru�����[H��22P^��{������6�a�WN8�L�u�E�>F5��o{�R~�Y\m�Ȕ.��K�Q�ց2.����/8��cG��B�+�%Y栠��'ޭ�--j��7��ml.���~j�n����©�kh�ؐ��=?�^J.W�Ս�8�"n�B,�U��,�qQ�0��'vI�?�֐`6^�fv����x�Bڻ�.8��9X\�7������T���Z��َ
��2&7�g&���:�A��˝�9"�&"6("����6�4Q���ܗ�^Q�Πn�V4n�w�<|% ʨ#�p׾�=���$�&����p���̅Uh��/ʨ6�+�]_� <�E��3�?���굶�&�Qg�إ�ɉb���8k�a�\I�q��V�	�؟mJ;�K�&��X���n
dn4���^6�~�I9���>�RP�3��NKb�Є�����s�,�ڪi��b�Ӎi�3��E�p� ' �7By����� ��Vh�cD�m���}�&�Tbd�#PE'����U���m��Ln~fj�~y��Sf�}u����C�Vt^��%nH�u���߁�O��#��D�B[�����饬����kTdTV�P�#�L�*I�S��x�:[��:�}r�9����0��Eh�ݜ(�t�� �ʂD$�1he�J��شЖ��P�Q�,��K�'�l��� w���Oȇ��p���K6y��sź��#���lp�E�����ɕp˗W���p�~����ަ���B�n�s#�w�L�.��0آ���I�?��������Bp�Nd��8Î�?�Y�k���%����?�����ʴ!\���r�c��������9��(E>C5&s�Y�Q]B���6��([�\���*#���D�Ԍz�yM ��X��}�&d;0��/�o�:rv�Q�*�o:�R�O����z��3�4���z����ٜ�r=5Z��_��#TILc�mK8F
��3��n��]r��d9����y?���1��$N#��Xpڱ�VV�$�#��A�y`���*)?ܓ��MHpu��*��3*_A"��}�B�d���RJg�>��s��p�U�?��3~s��"(��b�G�H�,�F4�	�z�iԱ쳵�1H:�jH��ڧ����W���ǁ�m�K�����%8�sý9�\��G+�t`l�R�d�׬��`O��~_<������x!���w�m���?1C:�ukC�x�I[.6dX�݀������Bb.`V�����3��Y0W���B���uit�������ORv�;�/��[����^Dp�.����L�O7�-�ei�Q��R����X����Ո{����R��̂�eE���z����=P��+^X�q}t�N�͞�+��'覨��uS'�Þ�9b���oؔZ�����$��W�MA�@
�	2f�"��6m�i�����3แy�XtQ3�����a�G���ӂ��
�ϔ�d���
��(w���R8G	���Y|���i��� ����d
`swD,��-��Y�Vr����1y_��~ަ�T��f{WPQ�۩!��������bf*{eI�4 �O�g0���y�S뺾�-�¿E�%N� �+�O��"H.�э7�uj�I1"�ו�2�\���硾�LV�����,U�0�*��5e�]6�ڽa}�[��� �ʲ��1b��Yc�=�����$Up���{5�Kd7·�,�ӄl�i�r�����Vn�7~ �F�$��� �p��U�D^�N7)�:��-���U�6l*~x��Q5��J�G��ze^{Xc\�����o���>��A�ʿI��F���)���w�Ξ��_�&:���9�������Zq0<�K�Lx�GY��}�|X�ZD���ڨ���	�*�^5<s��_8:��n���"���e8se���5gd�����AE&�'��jڙ7�U���J�H��̘����ӝ9U�ۗ}�r��}·H���I���Ȋ�f!��Op������N��y�YA�����?,�R� RR��h��@��<-"�&�2h�F�}i��r��`T��K���1�`L�v��{�M`����;�zk)�=(r��Mӗ ;;��F��aHk���Ң�z�Y���x҆j�ݪx;J�m7ֈh�d���F��IFQ�nҎ�-�C�<]H[��V7:�kJuǫ����}��L�d3�ݽc�X��;c��aX����m(B9.b��?��Ϣ�x���/ﱽ�N���ٮ�T+ޔ�V�©ƛ_�7_�=�WJ9�J�{D�M�I�����UO]2
��M�{N��h�Kt�v�H��P�[�!��X{�����^S��ށ�gnkR��#L�a��n2�����)V�ѩ������P8�>�oN����D~&���gnb���o��[��GJ����f���˭���e��P��"X�{d@�����Cu������|<d�O;��>��z�g��b���{͢G�B}�}�f����tP��}������'j)λ��4KY+�-��f��b"Dm�Q����E�~���Q� <N<��^�~=Eʇ��,)�׋�1�;� ���UB��i�Bx3N� Xqzŉ3�ͭRK�,���G�7�ʮ�f�rjR'X%�;��M�k�=R��_A�q��ɩ\e����)��^��L����C���O"P
�o�DZ(�+=���<�^�Tb��Y�o���V�M�A��ڂ #�;+�����c����"*�"�6[�?�]�I��CD�K �1��� �p��D;�
bS�ک��a��V'��s�`Zi�F��)���P_@_(����P2Y�;�)����С?H�O:�w�q10N��l_4Zuy��$2�\��6?�q5��$��#��֨ص'��꿊'<@�?j:?���A�&�$��Z�� 0�c]�v�ZY2Ӂ��Dm��f*=����������I���UA�x8�0u�;���6�[���|媁���xI���NqV��t!�J�N��Ks�I �ȏ�j%+p�G4��]�)�A�O��ޢ�hP�f`>���1�y����ƹ�F��z=.�h�G�����G�)��U��e�tJ�lT���ݦ��_3���R����t����:b��f���s
O ����x"�O�~*��S�����;"o���Z�����"�<�%�a���NQ����"��;��5�Ŷ䐰2˔���\P�N.��+�`�5'O���y��aY�/�	��x�w]|}���UW��8�e= ��]�+*x7���v^�Ƶ&��"sΥ��`-C��E�������/�e��KD����C����D<�	��3�S� ���lHާ��_A���E�l����̲���Z�(,R���`��m�&��G�G�圉yv��!N5�e�����\ok��Nh57���������~�QmFX���}�ק�oR��0�ҝ�Ul��k����=h���h�uo����+f�������N��>��nE޽`��������a��x�鱪F��_Zdoi�=�|k].�cw�0��䶇���mg�h:�W�J82��Z\����B�CG7�!�s��(�3��SYV�Ғ֘H]�<n��ib~��O���?%�-e���E�@~�V�޷�`x����P6oX�r�7���?ʤ3��%������:�Q��a����s���HW�6�:��,�^��7�^g�`d�"�S���0�W�}�0]�=��Y0���/-"k��Z���{xwRl\��!�~֛uiV>-�q��K$��+~+�ɡ�-��y={Wh���k&T{�k��룠��k�8��T�_]67"�Y���I����*]����0w�c��=�j7�R��)���*����2'��BT��(Ð���A�=������J�#��Թ�ʿ��4�!;�䙦��J�j�,�o������2�5��%m�&X �s����쒹w�%]7�zi>�z�HH]�;�S7�n�J��s-��X���>��<�*�y��v�b	�O�Rz�
�mJ<�sF8��-ݼ7+Z!��@�R�V�e
4�2GFJABۃ��υE�8lD���j����(8��h��3X�J� �3��M�y�p$Hm��~��7�݊�Ì>����z�r1�Ն��]~ ����.�yM�m�4~*������~q�����ͫ�j%cq���	��|s�@�Π��8������}c�}}�K�v�['	?�>#R�� ~z�t9ܛT�Ej�@�TP���zzCo��d�l�����]����c�Dd���t5�_=�)|�6�ʹly�mB����G�1r����筁�N�[�@���aR��W���n�2(�仠҉��ᕽ�wa��Z��pgj�*C��_?�=�4Hx�>���V?T�����U��5F����,O��ResA�_�6]��63��I��`�v�'�=X��p��	i�'��.Gz�ꮏb����!n�f�C˕��̎ʲ^��G=��H�Ü��K���'^��6T?4��',7?�9� gi@!��� +�4�;�Ʀ�z��o;.��:0ʕ\#��E(u<�M	J�d�^x[��x�5<��4H��C�S�Go���<�U��d\����T���=V�J��W��`ICE�V`0N����y�gɫJ�m�d$�Ϩ��õ3�$5{w-��7��4g	��R��.����P��KD&��'g�^�׉2^x��|�2��Tw��l:Q���}+�����S�ƈ���<A�H;�@�
�J����Q�z�}c�� ����i�<���@��9kc�Am
Ҫ��>���#��ܜ��R&��(2�EԢ2����h����l�%+'��D�D�ی��0��Σ�k?��kW�HY��rK���8p=�A����r,\����`D�YrB�p���u}L�B~�#�!���t�B��"�L(97=��s��ߨl�\����4�x gWE�[������;�^2	���co�����F��i0>ύ��t��͸k�j���χZɃ�Ѵ�g���Ehp:��>�Fs�ho`_P�D#q 焇L�*f���e"��-f� �p�M��Z(V:��A�)7�'���ò/~�K7T��GF����l�?2q�Hu]E�[���-��+���F��b�,�Č��y���͸ߣ�i�x~��}"P�X�F���ܱx_MD��V2��!������`�/n�zYVn;�8�-�% |BGk���g.��<��Rܟ[�4Ue�o�i�Qj��a5a�ü��)�@jE#�SjO)���f�J�Ϳ��ؘ̜͛� ١M8`za��	A{�H5PY٧+��i�v�6<L0m�%�(����Q��4����U!U����T�fu��Yغ��U��^i0��w�~����-�=az�m�{��(&��o�_iLxڼ���F�#���ʯawy[VD�F����@Z@{�6�hfDg��/h^d@:r�(�O�x,;��=Q 1���M�!�p�F�wi�w��$mM����{r�[9�z�!�Pk?�-���2-�*��@��KX�ĕb�?���t�e:��d�w��|ҩ��|�ɼW.�{.1��&���b�ꈒ+�<��)h�d�Y��h��.-F�^�w�����A
�@"��2�:e���nZ3�yO�C;ԿP�qw��3kT,�OҪX�a��|3ݷ�H)~IO�H��lgL
���^;V���;m��A���m��P���ic�,y,�yM)U���L$�Wy��a�q��#�����d���.D�'���A�%��ce�c]������.?߀��D����1f�vr;����M�c��4�V��43��
����&(����i;_��`7%q�Nue� ���x�>��3X-!�h����-b�7�����⛾�� �j������V� �<�)8�p˹�+�O!#�w�_I�KfB]J��ߪ�+*W7�4�*��t�M�Ȥ�a�{=B8�'j��a̹��jӝS�:
�A���r[�<	oQ�'�d�����L�IJa�(�#Q�� h���J�1r�y �p���E���bl���4���d��FN:"M���L�
v�{� Fq&��dvk���a����.��
bT�e�c�m
�0�ũ�S6��%]�o�N�B�bA��v�o��1&��j~*�������/)j��:(NUt�x�	)GYc�[�i����R`0�/��+q(�f����.��ҡ9 �h��]��
_���j�@���������N��ٗ����ȓ1Ѡ�����7��RADx��}w����i��M�<"D���Żh���P,�ɼ��M�k��%���<�
I?;S�����:J2L�pb7|��9��	��9\Z�G�z	N�!%;c [3BCoh��i��(���3�{������Ō��p�d���dmސ-����4 �D.� L�0���}��<�0��捆���>�s>�qX��� �2&.��=P����{]Ŝ�Cd"�ߣ���.Q��7DG|�����wϚ�jp9�e�E���gdհ���"��m�Y��M�i�}���r,Ǧ�����d�o����v>S��N'�s턦zf�������۝��Z�JO����c� q0�w�Y��"Ur,�l�'a�h������1%��E��j=J�`�K��4�m����h|ts�d5]W��c �u����:5*6�m��'*� ��-�{���KB�������KT�ֹV'�I�w[�����(Uaդ�)d�B�����Bc���ҐGn3��C��M*`'�Z�O�/s�"��9��a�i���̭�}��ᅉf��{4�@B��� ��^�PS����G}g;����v��Q�c��HRO�B_�j�l�d��^���l��=?�h���)�����d3���oم�|V֪�D@��r-���a��S�����u�����B��4ۮ����sW�f+��I�A�K�k��q䒟�� %�EAfIΌ�Ӱy��Gz��ֈ�k���{x2�F������2�O�2.o�ܡ����NQ<�t����,}?#�5���6^�v
�)��n� m5�Y����s�c@�f��%ne��w<��`1��y��p��V����Z4!����a�s��b
�uT��*'�����0�䟂����c��Bc�@A&9���Z�[vC�$Z6(�z���ą(W&��C����\�zXȞ�6��?@�T��[���7��8 ��T$�eQ��x�7��M��Gf-��5�riu�獓�&#+Tf|)d!H�O'ݥ��#�~�Nİ��Hvsm���g�zd��$�"f	�Up �b�B�
��Ϝ�,�-�M[�a�Y%���q���	4B_C���KHln`�H��(u�3X�	Ј�����[�d��W&q%�U�E"}s����<�B��>Z�o<��0��n�������rl9��,i�H������jZ�]���ɸ������ｂ��@�9��m���W�� ��&���ƚ�Ԏ�^(�)��+s���K��K�35����|r���X������*�l�<�Rr�0/�ی�Q�%�t ��5��M9��E���Z�^���d��v@�i	Q�-�ߍ����l�$9��-Lͥ���^�0�ԍ�Dz!X���ˡD�?�0��e���RP\����� $�\��_�������$���zu,R�1�{�6����"�u
�	y#�E��O��ő��C���H����nH׿OL��W�q����� �����A�j��nǖ,��S��;�)xB��ή�=�\��-�j<�(�7�;�1��O�_S��BS���2�*�����,ra����R;D�D�!vf��v'U�]��9u�:�Ӳ��ҿ���537����� �y��\��J�-_����B3y��54�u�:�g��)����:��	Y��o3RKe��<.$ʴW>M�����!BRƖrKz��KS�����$-�w�vtP��CV,o�`�g�%���γRԫ
?3%e�m�h�?NA	*����K�V�ȏ-�,g�5�F���A�^/��m���I��|�ÁE�I�� �q���x�Ḙ����F_�0yc��}4�a{�h9��ė��ļNd���T��~�ّ0����5h�~ğqҎ+z�<P�m֋
/��u�dw�����.1��a��6��?Tl���gu+�4����&S�MtT���g�(����� B�C��1�B�	���
tvj:�N��E������b�hyXpE�&{�k��1�`ߌ}����@l�3� �ߦ��h��X8�5�C���hiG.A�,(�׎+q$WO���ǂ���a�@g�5N�e��x��Pz}ؖ6z��$���y\VN��I}=&�K�v��̔����d;�5�F�~�tE�J�xH������A��]�Z�..?��>�]���Ļ���N^�ԑ�� ��Bj�b5�1a��sȪ����ڍݴ����M��c��5ʷ�Bv#_|P�b��������J�����	�~���%6�H�ļ�C!k^��v�������V��AU3��՝|�F)�D�>IbS.$��v��\�C`��fT�
3�y2!��j&�"������G�BF�^���Gt^9m���#!F����C��J%�2in9\=�	$˞9n�d��⧁I8���aK&y�M�$��8�z�� �m�&2���|����>���Y%�.�g�%��,P��;O{;j���ia@L���O�b��n�<hD���*��$��W�Un�z��'ԝ-��9=��}�u6~��"�ؼk���C�2L�`L�%ظ����Q�F)]a���[��\W�Vdg���3te�:b�1���)���~�θ��7U��y\�K�����{-����`-��4�ulEлc?]:��b@Z�"*=2�< vZ8E�㾽�ϾRį9
v�bꎜ�j� ]�v�1ڶI��$�!ª,~#�A�4�|!4i��V��} 2"<C^��N�Z'���-�N��iпY��[�e'��U��LDұؽN��u����r&2��R{��abq�n��y�������}~��iJܩ�6��K%�Rp�U-������p$AV�V�:�q�݃���>*���*�a
�?���X�U��i���U��p>��D��F �Ѫ�g��A
$u{-mR�7��Y��9��"�LG��V�6��!o��#�t��H�>= ���� �C�(�1>�aW�k/�e!9|󔇵�~%��?{%A����~�'}�״y^��%s�Sm�>���	<��E��K�>�s9lY-j�9�F�!Z-�n�wX��~j@����C�A�@/��l�C/i��88�<ں?j�(�-m$䃲��+u�O��m���ϊ�p��I�>B7/�1�[<��&�&=Q��!�I�mdh�Fm��p%����8Q�G2S�`U>m]�.B"M���?��-^[ �WQ��CA�]�ͻ��D0��)\ 3|DBI(�������ə�cy��Ռ\�K�l��d�{0g�����w��
�[����B���z�,x�������G�����Q��ј��e�e��m�ԭ�am�6��������|�LO��H�䩮H�k��ʗ�s���ͮ��лq�� :I�Z�gO��ů���S~���|��2$��]�*a2���klۚ��R�|�����T�����+�ų�z̆!-����;^�ML>MY�/��!]��m�Ma*e3h�LI�t�n]�2�l�)^P�yA���Q��Gr�v�y&���-x�q�!E�H�焁VvY���k��n��q�t\H�*�H^C�o�����Dh�F����7M���H�{r�	���V�� �ă���;^�W�&&#ʔ>0׊�F�W�~�g/�na���� ׌�ͼ);[��/bH��H7�B��"1�ptL?9c�0W��8h��
2�I'fB���s�w�/\p�4�ySwJ���Y�U'�&��S���F�5-�x����Ym|�B����e��K�vq��Ҹ�8��a�tQj2n� �t���%Iy�;���
�؇u����C��������}���f�/	Ȏx�kn�mE5"��ޑS�B�����R�N�k�Y��rcLWV}~���$}i��� �_תm�+�Ћ���=�ݦ��MC(x��� ��N5V<N�O�b[Et��_�ps�'^_9*�N�E'a�ʒ�y�TDS���� �J1��Q�7������@��g�!�o��̲ߌs���L��l�1�����(R���.��߷
c����1�ɓRQ ��)�~]�;p�[LS(bߝpg�/]�g��*�ZgA<�7��?y�������[o٠d�W�~�{�'�h&w�����X�ul�>�t@�QȒ�R"F���� H�U�"N圅�F�v�*��҇�W&�����g��3,A���`�KM�����^����I���0񐸨�::W_̴��ԭ�"Ʊ7t�pkV]����q�w��3gm�=4{�[�D��n��:,8�,8h�������伹�J[,��%��'��*��|Ў�Q'kU?�XDL�Q�vH�肎E�n�%ƥ��z `�Q�3���x�}������Ti�vېv�IІ�zs�_�f�k�t�2F42Ϫ�:9B�ͭ���P����J����!��lY&tq���$�=�;�WE��q?�t+��|��(~�\�;S���+�$B|g�eiT�J�#tg��"��p9��0�~-����&��C/b�V���Y �2�����G�&N��Y?Ye��� � Y��{;F��{'�͙[���B������:Y7�%�i��t�X���������u����fnGf(�t*t5I9��|���?�x�r��Akq��. AQo�t��a� �Vu�\��3�D�V4jD�>���,����~K���FK%��&�yH�;�}���"��i��&{(�����Y=D��o��m�yr�d��Gr�������k4�UR-�����Y�o�>fq��Q�f��R��k��
m�	3����L�\�n�[9�w{.y!�z�A������I�Ǉ����]��m��+�x駱,Yn8�)V9p�⬛�iI���,��a�5�s����֍�x�Y
x`dg�n]H�h�������E!�wQ��lҪv2��݀���]�52� �/��L�QO�oown�n@���" ]n)�'�q�x2�xy0��P�z������E�ӜdWZ�����C�g��)�B��"��z-��++�z�)Eh�j2O�Uk���������+ct�Ϣ܎��s��]t��oO��p��N9�a�k��"97����L�QnoLU�2��9J��S�L;e�1e�����h����x�nP�\Ł+���X�I}�>�n�Ё?⸆���
��`�ܷo{!��j��h���e�9���?���x	�����x
�a���K;3V\MX��G}��&9ެ��y^�$R��~Ǌ�p�q~Ӑ9 (5�v�9GK��4��.Rk(����d.0�Vɞl�������}�2`�V�$��k��QRW��t����K]6����T�diQ�r�G��"J����L*�>�$�b�"w�}�L7/Y8�N{�����"���f��O��7">�a�n����eQ0�U2?ר���v(�;xci�Ҧ���0ސ���H��+Z]��[zs}�����V�1d��;dYy�z���Å�k���d���a���l)�|"�s
���~
���Yy�G�R`u�i6�/�ucҝ��"�ͱ��?��
PqT����Y���{���]�J�`9��8F֑{xzu��!}c�_Y�\�9�'EI�K�.�xV�Y�ND����{��++�j���-3.�
14D�sp����Z����)V�;��ۺ�ٮ�,y��4�@���"��kV��^9�܁�{���e���9cFM����m_f�}���E-�(�F+�HMGV��	ׇ
��J�f����M#�uBS����Նl��uz����|�o�JQ�)��W���aG��G�5�S�ܣ�?�|d�\�v�£@�y�>&��2s��'C�n92�tA\A����BEr�u���m���q��d93�x۰�r�ߥ�����T�����I\.��+�w,%QqC���'z����SA��L^*f�񶹻��$���ZeTbj���<���qt�_���L',����ޔ!}=F�ߟ<%3�ίX�8$j�͟R����rE�K��4~�e�_��NzɽR���1v-)��g�u���ѠQ�� �c�'�oYa`#g
`��'Yjbh�Hi�f�>7,N��?�����OB�
�ҁ {�+�$g��p���G.���wКcc-S�}}F8'Lb!7^2�q��ڦ�:ǟ-����*Yu��yEw�G�)��-w:�!ػ!F)(V������M���V5���g&l��u'��Y-�ŀ��D���h�]��Q_v ���XZX�O*�G�����sUËC��|X�Q�0^���z�L����B��C�8u�0�h�L�I4i0��J-^�7�H����껺 ��N�uCN:�dl�lQ?��AP��GkP�����	a�,Ө��z��6����[�b��e�E��-�0�Ɲ�Ѭi����s�9�A�?��Nw�2w�oA��Q�ZY��l���C���~ ���ɲ�T3���k��N+(������Gc���]-:zdʯ#��b�������9�3�}��eE�k;�F ^�M������j����`-���Ve.B6�O��RONw�\.�LH'׉���y�����jT��q7!��]�o��d�d3����.W�5�1��:�U;}�#E��:��a�à1�Fd%8������,���;LMme�6DԷn&�C��P�+��4Ɛ.�V|tN:���`s��f�<*�P,���ʢ�'hl��Z���� ��s�Z��VO��IBZ�s���h��
�Џ)7llu<^e�y�+	��lu~b/��R��\7��+���Ul�S��B_m�<�;(���x;�B�z^P���͢��x1ށ>���@T��~��ȱK?(�G�˰���ա�[���Y �
P�������%SO�O6V����PP�DS/@��=�����sV�l"��]�D|�N}�VZ�/��x+g{Qu'e�ԞwX��*~�)�4!mo���%��1�݈��;֐8�?�[��cF��E|��=�n'�8���7����4�(F��,�wʔ��rD�ȩ2{��:���K�ֈ�x�o������18�R\xM6�+����0l�]:9J���[���
R�X��^��=�K� ��:�����d*Cw��~����R���c5EG!m�
�A�1S~8��h����Y�i`���Fi?�=�}?��W�v\w�a���9�*^*����[�و����f|���Ffz#�����B~�ra���
�p+�yT�0���	�Z� ��D�@���:�X�2�H��U�"��_��F���n\�T%
�63�i��c�8u�aRO*�����RAYl�eSKW/���T
����*�wQ��#Ƕ��bIql2�I+]-�xA&�_b!C�aj�����ԉ�򢘓�;�GUc�o���x������f�j�a�G=z��(lwLq2w�N�̆tݿ}mZ�4��5q�HM0��f�&��.�$�%�m��>�����s�B>�ɿ�k��X�Z,S��G� ��UPc���fS��ޱ��+����3���7��t�]el�N�eNU�w�0b�"�k6�3Լ�8hW��~/�'3�BY�E�J`��
�*ީ�h�\��<x����t�\]��d� �ؽ�6%"�\��Ҳ�^��3�\�B�~�PlX�a܀LoQ���}���k��ڙ6����3Pl�K0�9�/0���Ş`�o�eGJL<��z���i�f�:D@�b�詗 -�9?}Vi���_S�`4y.�k��JvP���,i*Vo#P���Ĩ>�FM�x��p�W�:�1�[���Q�tcz��N���F����(���]���=H�	�ýU0n���ɫ����p!��^{a�utw���! Bk����(.Sۑy�6�O����0Q�X֐�_u���r(&�����cɖU�VgЈ��f��O�]�`������\�z�z�^�2Og9@�"~�&}Q�n�.eʫTWc'��V2^���I�C��<�0Έ���z(��3��81:8�OVJy07�ޜD(�7*���zXن�oཐ���}��IK�f�	i�M�]C����4���n����k��|�a�:h8���#�<l���m�6ɩ�G�JG�CF�4���U�Q��Ř����߯Tr�%%�ֽ�"c��{3p����C��"� ���|�u����|$/�֙����w�9R�߬*���h��;/�J�k[%]%�:,�l ���kC���������1hc:��Xq�����n�	:�	#(A?���h����u�]�E|���N�2@J�p�vg.���Wc�JͥbЀf��#�����ʦ���c�L�}��ZYg�������.±rru~�s���dgM��:h���{�����b�%��Z,��/��RW.�����}a~w7J�Ӵ,6�f&4��^���\ҝI�pи��(0z����{HB�By�` v���O�3L/�"�{�pH��a�zp�*�
sos �A(�P}�8^#�~W�24��P�scި���9����SCm����î���?��(Q�2��y�6K�/�������;,����DƐ�p���z�4@�I�EQ{.n�Rl7D*�9\�������xF'�y�W��U�&���yK����\�(��&���2��8 j�l���@�!{&e^�+!6�Zp����Q��HU��.?����:�F1�@��ޱ���A���ՏW-B�4$Gp��*S��pvw�ƈ�@7��Qx[�o�h�ڗ��i�[Ƨod����4�l�{�<R�_�i��[��>`���x����Oc�s
RP��[c��8����ic����	�����	ҞJʈ��ں�rB�f��`}���͙D__�rDF7�	�Ա5��ܵ@h��v;<�;�a��ԥI����\��k�`
P��.#{��=V�wW��EE��
*������,���J#`K�/�43�dU�������]睑y��r�,v&�����߹�δC��+KQPC�:q_=��b��q����+��|$jI��O!�I_�!b�'����(�����~� u�ܸ�[.��L��p�I#^��r���Rd�8�g�p�s���E���4<mN��q[�l-�"�l�F�C���C)�h��8o�*���� ��]�m�[�K>��z�d��\�r 9+{b�r|d����sq�%f�}���t{og%��N܅�v����꼐���;�e�'2*����ki=�r���J@Y�Ċ�=s���g����wu�-�����1�z�G·i~�zf���Uچ����yk�d�!�#|3FaMI]�c��.���8�t�w�ӂ!Y&�=��^�� �g�X�p���P@���yxx5��kQ����lQb)�n_%�P��u� pYZj�No� ل��ȍ�/!�HW#m�zWl�$���"�N�Y�Y3�.�Ƀk�������$��j7Eo���sA�&+X��f�g�<�7YK�k��@4�j���+����(�I��βp����y���+b�VԘ��CGն�Vu�R%��|�:���J0I]'�X�L���4�v�p�yb�m�"�*�Q$��g�L�kH�g�n����^F���6��^�j���d��3�%aE�Rb(�
c�40bp���8��6�9^C����l�h���-��c#�k���_bC�A�y󍆾ߝ�,��f��=M��η�!�h��L�1���iB$RGD:*�����&`��, aB.�܍������L����3&����*�8�e��_i^����0��9���Һ��"��X���Z�M����F��ǣ��t��!�c�c�o�y���*56�����V�1�������#S���(���9��8*=?��FwQt�[Quc|��0�/��L�84�w�����^P)R� ��T��_�Ї�S�����T��y�f?�7u+���!�X�wW�*ZeE*X�RU��y
��f��8�C� U���ՒÔ}�2��0 �KU-�:�U�����#4��d��`9�t 6b����"3ef�0YJ�1n�y3�,g�i{OL��,��~�� h5������)[�N��@��1g��'ޏ�|y:YvK_^ ����c�!�8�����Q�����\��T�-&�A���}�ծ d��>L3KN$�9��4 I��Է-�i��,!�W�9�Ԯ^f��孉P��P}0�F����~r8ѱr�LR����M��37�[f#�m�#�g��N]~y���\�Tɜ��|��eeJ6z���P��.���BB��0��j�h�s$Cñ4��p6�y̕�������өk%�UOe�w�'6;WJ�ى�%��p��Ĩ��F�O,'��z�J���뻲�p�|
"
�{z��f�T%�	6~�j3�|!�Iz^�F�R>߄Z���+�,��Z���b���{>Ҽ�(���QԔCd��S�x���Tɱ��H��	!�8$* G��{�t�ki[��0��H��~~� ��T��o6S*ǧ�&��Ѣ��{�d�,f~����eP������+�}`a��B��$]��.d"��%	��"p�'{[�������ꜥ~ܾ6i�kG6Y������VbX�{���]�)�b#nM<Z\@���M�����D@��u�0�~�8�K�1��H��C`����yV���\��������͟�c���Q-���T�p84`
^q��dRH�K�';Zy;K֕ť�g�q���Ys��9�r�Q:9�i�=�ga�)ԅ�:~�l�oRj�d�8����﮼֛��-[�%��~4�6W	���"�4*좙(�G�k'��B-�-�	�I+�,�8S�C��,����$�:���8�^C�!n���M�����]���_��p��x�%o���R�V��l��5��\�q���H�,��7�q5-��:QS��h�V�PLjR:=e�xb3w^Dm���ٸ�My#������(�ֳQ��z�\;��<*�=��tBHKy{����{r0MMI^�F�#�:x"�����|x��|�þ���I*�I��4�c|�9}Ľ��G~�W}�tD0%�:^n�"���%��U]�}�{"���gz��V�T����l�m �Dz�j^� ��y:��>0����=�k�]+�x�Sm�/�d������HK1�z��E�u=�I�Yx�mw�տ��sx�w2+�Y>����P�Z���V*��#������	�Ku��3C�3+�1l���tH#�{&,72&����ǿ��
;�E�z��	�����?��x�I|GN�߳�y�z8x#�J�)��g\���a ��Vl�,�H�s��B��X����=u���Մi���i�.:��vY���lp��`l�Mk�� � y�eH�q���T��� ̓R��-�4Y4du� �+�1�Ţ�R�����;�6���D�.�H�,|�toIhũx�zw@0�<�I�!S��R�qq1�6��y�gV��@	�!(]l<oQⷝf�i4hD�9��w�3�V�l��M�J�Sg�6E�7�alģ���1��'�����X�5kiBߦ��7�o�rCs̰zͰ�t�Κ<X�����X�CB�������ߒp� �Y����% ��o[pE_��>�'+D�>g���A!�k=ҵ�pƉ��蟰�b�U���p%��~V�w&~$�s.aj\�ͥX4L����R��3�Z�틓�����&h�8�x � 	X��ד	�AOhp�>��W|�i�J�u[t`�i;Z�b͘'Q��w�)�I�?���W�j�Q� /0����B�h�"�ʧOm��`S���6�ڦ!���J1f�0W3�A'� ��`�͒FN$Q��~-V�[nAw:G�������2;��Ȉ�(�'�_����ڭZ�� �R��H�������G^C����@�+�gѾ�F�a�#W+�.:�4eI�L ��jU
��8Zo��Wa�p�Y�D�����Z�!�m.���Q��#ct8�_����:�I��]@�l��N]7��{;kK�5��+���W{�]���\m�}}y �@��_ �7R��0���RC��݊�l9�㬜�~�������w�e��P�;�{:P8*_GW ���&PO�q#��&�1+���o�E�z%"%�7�0W�_n�d�%�7u���I>FjTI�з���$,S�GL��Y<W=B�:�Nku����cU�ȃ�1��䬁�ZdyT�Ħi��e/�ps7�Jʺ�&��3��$��<����_+za�������m��ni�{�(���i?Q�*�G��W���Z�t}'��E| �v���-�,�9.}��<f[Q��λ]g�e�<�1[USo����q��T��R�.5wj8��0��ف��p��Y
���z�f%��u�F�؃m��?�y�B���L$cyr�P.Ǻ�2Қ���8/]�s��À��Ү�����>����tYւ	�1�V��G��h<&�-#���Ch�Z�����O�7��B��*]'G��i�21�J˝���I��< ���}\}��r>F�#L�_��o�qd����u�W�9��8!u"L��F_��40+������a�PG�ة�K-1_H��O��?"r@�0���tSNa�� ���l�1���B%"��φQ�㰇��c1Lb��F�'�@KM]�@�ԫ<eg�u��9X��[2��qʷS6�D���i�-�Hr��)�����"��Tǜ����ȡ� k�b�� ̅��rʦ��*>�x�r?��4_�o��$V0��t �V��Ez�1����Xd̂J��:xG�֥!r��L�����m�n�"���&���RXK]C�ɱ�� �^zݾG�$��|Y��0(��J��QYЊ��e1���Ê'�xS=�_$���43�,6ݒx���A�ߢX��
b�ن���[�["»�B����U��Ƿ���3���$�c��$�<��yFߍ�������/Tl�nլ(��#͐_���rT�a[���nA�����EJsˮ��=C���L�^�C1-;n���" �ݪQO���a�2;���l(��ף"^����05A��K�Rg-������u�-����� �/k����(���o���yv��S�UY��#��i���+\�SX�,�ZL�n�+#&���'e�% � ��yZ��~��۴MgNYv;�#���:��:�,f?�<O��dZMY~���^�ݼ0"vm���ٝԼ pn;����D�� ���s��9�%[���zP��<�	ڼ]0Dض	���w�=Rk;�o��Ph!/!��vT�ϧ�
���]"Kf��;�c�X��s?�a��hdZj��
(�Y�ݔ�FO�`\�P�UU,%`Y%M�.����Z���˽�2f���C���̂�;B��"#�! �1I�E5�zo)����k,�U�l��3н{R{N�ǔ؇�_����b܀��]�F����ȕ�i���a΄�ڎ3p�b����C�0	�����`��g��c{���f;.�5�Z#|,c�2��'�|��X�_�*��|r`FR�+3���? ��.HR�}�EEw���`�:���r�ɧ5����M0�)T����أ4�ϣ�jI��5��lr��D�k�ʵ`g�:����-��{>لNRc6�/�XQ�D~���R�V�,�2�mOU���tC�GUmA[�^r���8L>��f|}�"�>��OL���8̀NJ�X�q�T����@(�s2KH:oF<��Z��ș�Q?	�@�`V�N�&D�����ǹfʋqѬyhe�^[���7�G�1������
�#=$Z���MSQ%c�����]Ukav�)�E���5��o�6Zx+Րߧ��>ǀ�c�mY������!�3H�h�,�	�����e��\��.�4�R�����,X~eW����G��ၝ�Ts��)v�Ӽ�'��0r�(R>�,I�S�8���ġ�����n����w���EL]�����;�Y'�⢄�ॼ��R���N��ū����.uN�4~���_��3�ab��m���FVn� Jb^�@z�� �Lݛ�]�cD�~]��Au}���p[�	%Z�\������b����c#�:w�خ��ͧm�ư@��Ԁ�C�+K+ׁ��n}ÔdZw)��ΖU(�!i�<�k�P�52qhؐt��5'�^�x��n{bOӀ����h��	�"�R�"��aw�DK��f�p�;r�rus��,�߼���]�͖��-��{.q��t�(g>��%<�����6|�O���k���R�lȟ:p֒]����ݩ���� -�$E���ٔ�J(��1|t��%�Ⱥ������\Q�^�*�
4Ք���A��Sf�_��N �L�8.P�<�[�%���G�X�4�G�XYkU��0���NA�Q\��_��?Sc�Ic��X�`~��@�����)`C4�S0����6ؙ7�?��'�����'DJk �� Ն�|s�<���Mo��Ӓ�8��5�(.-]{����v����jE�`���+jr���O#b�ڇ���{��>L��|k��s���A���p�)�]�̗spbEU�B8QgI�$�����+i3��*E���SE���Q<������Ө�B~T��7ţ��&ѱ�}����t"�!�6 �$����ˇj�/ͅ�he���� [ݷ�/V��C�1P!21t��o��tw����%Hn�6��80���y������A��Q3�5E}��#�]��S2�}Ʋp�P K�2E�F��#���g��ǧR"����~
�����ڒ�6*���?��o$\`�qf�2����ZlRq��!+^v毇h�6�t��fhK�6FH����%�r9�{�w��=�&�$�����[R5�4��~�Ŏz�H��0B�Uq� ������b��[��L����s���䲗�����mⷥ�	�D�����b���rLg�'=�yM!���9"ٖHz��T��@��|>��m��Nn������p*��Ew��%l��dj�|���ŮBa�^�&];C�;��"W�=�[@d�f��Ϫ��"�q���~%�B�RHy:��E@݌��y���Krt��H$u%:=c��<G��o�%�n�{�n�!�	���b�M���w����G���Ð�mQ��f����Iq� ����$�E�����)C�#X�CH��R�im��I��x��҃���!��_�����=�Am����¦���P���(��8�oK�Z4��
�F`(Bz��V����ҵ�ب��yG�K^8��P�O�H���a+�X�
�Ym>�I_���p]��6q�������_�@o�����4J��o���Jd},����jԮ֯�2Iߵ�(��"�R6��1����|HR�����&]�2)0"�`WZʰ'��1�Uf"��,��t��d`b [`�;���>���#v��[9\S��x�y� a΄��8k��8�J-�
U)��$$[IN�p���np�a-##�-�-����Zu8�<(n�wbT�_��'3Ï��}=���u.lB��l?����f �ë�>��Jzh��R!���pH�@�5�bC�T���1�{y��͘�T�px4/Y=�գ�L�����l��[��㞖��O��SM�S��.Qͬʖ���m/[q�JzHa��Hpv'�����a�7l+dtp�x�R��Vq����U�#)T�#�{�w�e���֟���M��b�W��=�L֣��U\ļ�t,}�c,]c��f�m�rd`�#��u[���Bl��h,�n{��R�i����;R����1����e0�����9�]��Z���1�j��	,�[�jþ�ɳ����Ha�EJ��>/�������'�a��O]}MvW���ͿY�}{��2���|Uh�Q��L�I��㲽�JA۰h��*=2ˇ��	{����Hҩ?�ю��=��ܰ�����F�y��u�ǝ�V=���P!I׼O�8�)ߙ���w��]��gy�"��ں�H/{Z�`��Y�W�$�E��ɤ�O��ߞ���Ӂ��%��$���-(x���t�+똸�m�j Z���/��QQ��Ue���6�=}r5�y�X߱���ısӣ/�P/�Z鋚@���
�M[�#2X1�'p�I��m����d�j�f�Oר���dL;�#��\�Zɏ�g5z��hnx(�i�#��F�|Un<�2-��E}5?pw��|x�IM
L<7����J~�oc?�.Z�r$�R�a8��0����A�,���)�������)�U
�]��a�n���"��7b|�&S�(�.�8Z�	��c��o���+��1%�a��X���3w��㣢K¸�=�7�ݫ�>O^�c��#�E�qS��tO��~�������ĴS�7�"��Qx'!M�)"��D�kFޙ/��.A�?�-"���M2�0�{����cQ��;э́5׃D�eG�����2K5�"����v�`����T~�O���rbm�����������K�\GY��(�||*|{�φ�7y�7|&+ ����ѹ�4;S����k�� �-�W<Z��M�y�5;��ۮ���;�t�d=�GU��u�6������ �'��ʜ7q����:����t���XF'�Ʉ9ܯ�]�[��m���`BzĀ�.�E�H�[2�e��U�/foɟ�X�$��p�{���/���36}�9�x��{����.#=�#�18��y^2i%�Fuu� 2_���O|���Ahປ�!e�<�~m/T�U�qmj	Z��r.�N=��%%��9�-̡Dװ
���s��g��%eI��h��]���gS*�csO[+�� ��Gǋ[:�S�ph���F��]$<oqyK�'�I�y|��v����y�]90v�X�� �	��h[�hvq��^�};�>|��x��,)c�l��z�Y��u ���ڲoP�@�	��kɋ�p[R	�l�O,�h�Mo�jP�k�=>��`A}���h��:��՞δ|�[��V��ga�S�Y�Ò<��ڽp����������e��@��\<�z@e4�N��1�7wFޏ0;���í���U{=���g�j�/á`���9���N��I�h^paK��a*!�X݀��!�M�+U�c+�`C���t�g�ñ��J�&��5XA��u���j�3Y1��'@�Iޜ�zJ�$�WM������)�	9R��m��z�����,����
���ڢ��$�D��bݖ��]�uE�ȇ�D�3���0:�GC	Q��/_�&�x퐼�g&��h9O盘,�?�+�D�D�4��&H�"���;[t�98t�R	��;tu^�/O��T_�H��^*"x]o��G�b���@�ʨvam@M{�'}��{��鐲P�T�0�^{-�ʃ�z��V?@X���{֩���ε��M�/N	��Q����0�.xX,$0�\=��I��L���L���aA-�� ���h�D�?d����(�eFl�2<�]�o�S�7�=ܺ�LY}��	ֺBy����y�K�'b�H-H�aj��3>Q�o���z����C/ư�KSn� N�ͮ;E1���~7��;�\��)�������I���˼� D)٩J`i���̩��)5}w�u,�CtV۰h��3��sF���蒷�����Y^�~7 ���y���peb(��4ie�I�[n�Zx�ݺ�;��L�	����J�;�#W��5�H�4r֞.��Z�o����[��M�I�<7�����`�o��w�&���Ƚ�Q�.��g�X,+�R�A��[E��ݽ��!Y��NV@�{*�=qzz���Z�%(!�0P�$�oZ��ȹܴ٭�Je�s�%s��8�a/�G����7����<w��ػR3g�o�e4,UL;��-o��"�.���Q�1�xR�W��0�a����Hu�M����/_ݰ(�]].��
X#9 }b��~ș
��N�a�^�@��׆��ŕ���+o�v�w�NirԕW�i��J���f�V��x���1��pu�RAW�z�V�p
S9߀��� 7�:�$J�L����pDE׆����;�ނu�3kPQq��g�fp<}�X��*p
�'��8�oG�8�t���xL>�T�Mc�;������ˍ�{��}'�1*U±��7���^Ee��u���6c��� `Vd�mifx�#��7ya���+?.-w��M-��u�����dDdeO��b�O?f�l������i��u玊��ny���皪#]�'2[U�z|	l�*f��;u�,)wj�Bv ��M��׳!i�q�<(\KV�_]�[/wY�h���t�(�I�]I��f��JY�{���?��q��a��sÛ� ��i�RS,`��j����4� 唬YS�(��r�>jr"�O��X�Y����9v4#2:����v��}^*�<��y$������+����M*�eJ���5��h�V"x�W�cs��,ѥ�V�iz�"ULU��׺�jq��T�#0Y��JG�і�H�PW���L4��:<�\<x�-��˯�D��?�G�������!��u����- Dh�R/���Mj�9�-_Ft����Y��f�o���k]<_,hUfi7�k�&2�Y����SE�]�R�LT��4Ϧ�݀�ܷ�[l��hyL�����3i���%�`�S�'P��K�uR'�+i�%��D�Fw�fB ��1nՏ��&8<��N��6��D�;6��V���5�F�Z%xg���/v$S�2)m��?��l��bD�^c���v��ˣ��u �9?�/��t�ct7�]'#͍ݝf"��}�t}�=��n,o�LD�C.�Z�̋�y3��W� ��j��OY(�dI-ۏS�p�I�a�L�~���<\ߎe�whB��x�~g��Ɗ6����X��z��Cu�+��c�`�p���ׯi�Kb�(e�%?��7�*����3��v:]Tc�I�H؇�R�ӿa��19)J���k�f���`y�Zq7Tr9Bڟ�JG!���;9���~��\[W��*i�^̩b��(w7�]��W���j�W��<��O��;	=Pl��e��o�7J
ֈjC�9��ai}X���\��̩�ـ���`���������F(���7{_;Q�*�<����@1�ń�� (O��F ��Eg����~�a��tDA�Gid�s���}�j}�hXV������z�����w3%�MhoW֔�f8�7˧:�{-k���-��&�Z�!��G��U�(p�6�ǉ��d\f̏�&�	����e1�"Y��N$�?|_1OtRŕ9���kU>�"�|Q�Tmܑ'���d+uQ��Ӵ]�:�[�?����P�_�ۧ;��͟"��q�g,\����J�����/'���sq&���K����x�����n������z�cH]��壦�K��KJwڙ
O��l����s�"I��;�؀S�+u����@�\N�N�S����)���Q�}rv��x)эR>��x�nG��᫚����m��z1j�\Y�����0��l@�8(��~� �%�8x�` �cIP�i���T���Z�����o�� 4&#4Xb��W�V�JJp����* p��3}  c�.�G�gk�1�ã��i�i�˖���%BM��.i���%���	��f�Lv��ϳ-����W�.>H&'F���9m �A9݃,��ZS���O�d�`�����pD��ωz�� m��J�����\Ri]~���L�ۥ�Z�A�ھ8����,2&䣒݂�9nS=
�\),I%�A8=��ɏb��S���7�u�]��聧�ߓ����sە�P�6퐙��x��w����upx+1������ɸ��)~d;��U�X�H��>I ���p)Bμ���\z��H�#����,��1Kgg���H;��#؀9�u���ّ��\�����
�WښJ���.����ɠ�,��H#x���UT�]Z�p6����ʶ�a�̳��W]?t��3�*H��U;-y��(u���h���R0rT�/�Nz}KB��=O�����@��]_��Tur��['�/�&��iq�҆�%#0o��K�;��z��~Z!,6����~�p��Ul�խ�	�
�ln>�zj=����D+��6�<?���ۅ������ȉн�@�64=��y�{C��X�B�.`~W*[%����� |2����.��-�cu�q���c�l�����;p4mһ�Vp!ɥ�:��8,<w�E�uM���[0��5PŐQE��#�Eh2ɪ$-/3�������z�T�w%g���hυ���[y�?٦�����\�K��\��Z9|���f�N�����[�9�hh䢺/N�"4��:���!�X�m���R�/�V���џ�kFu	���3Q�l�`c��1:D���t׬���\��G.3I,RlMK4A�D��d/؂���H�dr\@Zt�v_���3�
ň������y5<ؾף��������teX�廜<���h�r���) ,�E7J�ſ�����F�Y�L^���}x<p��
�@���������e����yPk}�=����}o���?F��Kۥ��W!'j_h�UB�HjW�1���\�߃��k<�)�4�>�.��\��0�j�IOpE��ewt�X������t}�#�&��	̓�"y L��� pD�J�@�Kp�V��c�/�6I3���rxG��>��z���}<������v�^����NzN����?��e"��.��u��M��P���*4H�x!�f�H��̏L����
s�ڝ�z���^�T;�EŃ8�����4$ؤ�����=l,N{��!�y�
SK�[�t�m��
�?+�\]`h'/o5ͩ�ڼ#�^��2R��s����H���/{�:��a�l�8z��@~a�K�_oD��De��ѝ�3�/�I��,������f�I��j�#H=F�+�'�^eb� $��ԑ�!�usC������<v��>�c�6M���Օ��ݯ^��z�1������1������2U]��U��k`�[�o�X�,e%@�]=��a�9�	��5��_s�Lu.YF������|�Z:l���;�t��ڀ���`T��a�Ww�O�EQ�ye,7��
k.Dk�y1.3�U�sL�%�nF��FeT�ee�Hn�O�Z��8�G��6	I2J|���@��W�Y���~����^�7�
�^>��F!���(az�d�hn*��Q�j��*�c��)��Hi/��
�*O9���CUD_��'��[8����P�:�qu�����j
���4
�Tq��|��vb����πƤ��Zҍ�9cQ�qM�I����h��I�NH�	�f�T�&g�fs5o����Q
���xd�����;��"�\r��D@I7%�� �4�����$�PF�t����g���X�e чH~�4�T����u��E)����*�>!;�����!nP�]ˊ˻>��#T(󛘧'��rbD���Q��Ŏ6�[>�!L����$H�&���1x�`3it�s��@�{��V��i��������5�W56bU?ԫ��Wvt4��#U�|n�����)9̒�n����l9��VJ]`8�ys��Sѐ<ޖB8���l�q}�&�8�x��;48];JU�J�pQl��齛A7qx.	�6�x��Zc`��zY���!Ē��[��]��wpiܷ� �	T�i��'�G{��mq؁"#���P���$]�^ςM��6� �7�{��ɡХP��7[�	|L֏�ޕ
Lǅ����49\��7���	OҬi�#�u�5ź�hF�G�
�z�I?v�;�cb�h~�� R��@�H3 k��K��Fd�jc�Ǻ�qF�|�"A�i�f@��{�]w4C�\۳���9��׽+e�A�ȁ�__��?P�Ł�Y��ԓ�]��z� ��U�%���*�sb���Ā>O��]���$�=�׉^24�a��#?��7B�Yc�e�6�2S��ʀ(��G�/���%�h���E'G���dn�\�?
�d��ϕ�بc�K�w֮G]��]�ʂ�Z�E�;v�? ^t���N@n3�}yT�&&���^� �iE���:՛��ҋ9��4�6ú��LQ.��z��ݷ����	��"�RsTZE���bɒޜ0�R0Z����{;�S������!�tj�;��*�(�2�r16�F{pQpߍn+Q/UZ=���m"�!��k_4�S�_�P͗ǙG�'<�ـ��R=�L���{��W�I<'7~�
�W�o~�Ҙ=�*��}��9d�m��1$.�YW2	������3	B����9�/.���9~�y=�U�f���v�f�E�+J;k���Z�n)֞�!4���c`]�(�`����$���+�l�B�"����Q�[v�e�[ܩ��/��z�w�$(0@�5��m%R5�ٚ^�M� �%��m�D`|��ˏnq�!t��k������GE�Հ��7tF�eL��Q���J������X�ܺˬB�Z׺]��j�Η��~O�䆯��^W����h'�
]�~&�N&M��j[JE<�GՄ�(1����L�inz,BM����vuy`��J�}���'�A�f��q�M6M��Ks�az�F��~���7�-������ܸ��ԸtJ�j,�	|}�����.�����Pw��J�pJ:��B�_��f(TF��=��_�:Q kA�n������t�c8��C���D�g@ur��K���[��^2��b�
�堛�v�b_1k����;�c!���O�*Z�i'��s˔�X���_C����O�$؞t�İ�����Ch�֎�=�p�s���3�s�t�L���� �}��1�CNۿ�.P`������#���ݣܼF���Cy[�҃=�,4�7z�Z�;: g�ň��'�e(��)z�/���� �]�֮Q(��oo߹�ۥ+��.d�,[���}���e���#�k�ЎV����o$7D��OGd�6���N[�3�	���U��N��QG��f�F B�-��Ωl�mب��ŷ�T�O		6<q��:�(���k�h�����q��~����>b�|���z�	n���q�ŕz�5J���W�B�9��QV����P_��_���ՅH�4�����۬��zV/|���Kŷ쿪�<��0k��$�c������Ҧ2��]TZ�A�tK��{�_6�o+�u�3��]Ja���$�C��xL9?�#q�G���K�dL�
��z� �o�����ƴ�Av\�`0�5�8�2��c���OA(,]�*��S�FTL���Bh�F��$�٩�'��ܠ�bB5M�Fճ/�v�Do������Ьm�@l��>pÛ�a�b�����5��b̠�`�h�7,a� �Z����<�J��V�6��X��������ù[�dY�Fo���H�o�h*ZL|�$ޙ~nRN/|[�\��2󝄤�$�J���1�#'�KZq�l��Se�7�����S�kxO���iu"`r��ťH���}� ����T�Q�{#Y] ��8��U�ŏᑓc���9�Ҝ��Y�y�su���p�H�{$"	���"�QoB���J�����)���6�1�Iȥ����$�t*�^�gې��s�>� }g�q��Q�d��Ԭɀmj65^c�vkH�n��3��$(yrX��P+SPZIɐ�P���w�N�#Gb�_��r�Q�w*\[���5[�N�N�\=�87��\�r#W)�h��%�P��b��א՞N�n&ҵ� �{��(��N������zD4}�y #MAe�m>#�bo\����=Ӱ�6,���w���
6��c�#s��5��.a�!���+�^S��o��M�Y�� ���h�?�:���6��\�RKa��9�O���2�p#�i��6uUݭ6��`��_4�`a��J`6��d\�ܹ^��Ȟ1U� ��8>[�jRl0���=Z;��Z���Ɉnyx�[4K�,���M��ζ�f.s	�%�e2���>�kb����l,��w;�����[)���-�'�o�vǒ@+Cw�"�!Hx�"����u�)�dH���+��U�_)%%�'��*�0.�P�n�ox/1�M���d/u)@�G�L3%���+MZ��UQ43!{ww����g���0$EO�}����Hh��V�怅�Ô��MxV��8��w���\����� ��n'��8�Ԟ�D� k�<�����7�:�jA)W<D�;�˽�l�4�MG�~��84VA��.O'�@C�1��}i�x�.�k�	9v7@M����KU��sZ�<��DM���>��q����*���6W|R�$��\��7�(��~��Z,�?O�bݵ���2�XQ��Q�����!9_^���فF:2�MpU����E��yu}�\�L^вz;A�]ɰ{^X]b5�кv���lc�]Aƪ��zOE������I���l����y��"�C{���)��̈�����������y��T�MG��9�MF3���F�Wh��
��X�k'���D���ŠUZ�]�Έ����C�xm6�sj��m՘���>(w���ޅ0o.*ؠ��K]U�'�CtE�'����FnU���TOE����&g`@%�f�q��ڰ�d��1�>�i_�ė�ܰz�f��j^�b�{Ĳ�����=��La�w\���V �Ԧ��j|�QFq�`��HO��X��uaڬ�r���Z2"R�h=_�*�g�.0�>��|�S�/z������w\[d6�09�څ��0�V����Q%]	M�.�>�¨!K�DPǁ��̪)J^�(��aK�����K�~q!�
�5����=X��SUr,�*@MLq�eS���a�GZ����72n��)ņ���[���I�E3e�WYLmU2aZ"�Ԃ�S��|��Ƒ{�ΒF�5�����\�<c�u�������4���:IR	"S8�� Z�{��4\B�^����C|z���2"�$�1��ۯ���<�L����"-���&H� N:����/�4�T�F_lg0�ʱl���ݢ�X �n���Ll�K����Y���MP��߉��Dw�N��k���l,�v�|�}ƣ�`Up�;D]�ϗ��{DID^L��8��S��f`*��n�����/��*sa��n�c'+�I�����L����]@k˛�"��/��4J�[m����I��Z�����٣E3<��v��5t����,�Cl�å[��1�ֱ�>FZ�2dShh���yT� )��M�e Z�R�f�ݘ������<,Gt���3j�y�%V*	������D�\w>�A:�k�����$��9e���Q����v:�"�dQ:Fȯ>����ރ2��:�Y��٢�x�z�l��˦\z[2W@O��Y�$oj�oz���~�WM#��6�
�r>)��Ŋ���=%)���c��Ϲ���.k��|gi`�˴x�0z�w)���D�6̕$۞t���>�i�"v��"I^�������w[G��ύ.��Ln��Z.si�;n�vb$����Y9�?��c\�	�����HkV�D��A$�%���mX��0�+��5w�����H\��*9�q!�ʃ�O}����D���MJ��}�+�k���D��<ݺ;�B�ՙ��#�����M�Z�7��o�i��Y�4��`�SC��0���A�����J�-�aP'������v�����<ؖ��_'����<�7q���� �V �T桸���f;�8��|�'@����0�n4n�9�%�IA��&�O�0�W7m��)v�5�`�JBsi9���ՆH�ť�x#;�q��J���[� z+�Q�k�T��Y*̹h�+��9���?��msv���?1�(Z�x��kL7��
0�"����}zd�2X�m]_�S;L�
a�^0&/�΍�</o�Sfo�ޅC�O��aQ���2����9��Ot��X��7�`�	:� <g�qx�CP�N�S�^M麞��za���-���\P@�����~�;�g��}Jw�=/,��]�Z�;��!�A����k`�H�g�����&�Vܫ#��V���T�eA��P�����3s�?��/^���Д�A�<W?�/[���x�G�D�����/T}�ھ~��q̪���l2�-���Y��@�MG�9R�x�"�MD�����s�ug(վ�W�ʣe/M��x�I�y#��at<�Z�����m-]�\<"�x�� �jj�����,y�L�Dۣ�T���r���:_
�q��A7�����r��`�!�Ur�<�[ԃ;6W��~`hsW�������]�� N�y׍�1e{(���?�R�A5��Ӫ���O�Q���}$l����Xo��b(��9�a��̭�i{�oٰ'oTT�ubio&7̵^�{u܄�e0�磂�=�l���-�I0V�J�I�d/�A= �I� �bt6
�ߵsS%����gtc��5j^|����!��<�U!?�KИ�5C�X��F���zDG�-�t���^�߼f�!ح�+
��>u$�{����o���\ӹ��\@����5����7�ui�k�Y��CnwG���/��&D��
,# �*���ϡ�|������4�1��#C7�C�e}K�fV�*������e[db��6şbp�O	��Os�|�C+�^̼�M��x�+a�Q%�x�f�V\ּ�N�*���UPUe|L�Q��S��]b�e̋�9�+�A���)�Q�4�Q��3�B��=�9%���0ϋG�G3|�0��r�-��߹z��@h��c�8bl�#q��2i�b'UCK*�܀l~�,���gk]Xjp�s�օI�� n��\�*�A����l7��B֖5�	@Jg勒�ڔ���/�J1�K�mɔ��	?��Dc��?��N���w��e���E�K20�e)+��'ö�˧t^vٖ�C�T(��� �K�Q56��v�"^Xd%d_�	�!L��G!��O �ڵ/ �)�uAP=�����7�)�+,]aA8	{��9ֆ�}�7�slw؍����%�L�,�Ň�`�`�`w]������iʆ:Sm2ئ�TG��{����u
���D�㔽W�}꩸�x@8��&L,-�\ۆ�\�9gE5�ۤ���֎���K��Ip5�"l�0���N��S�$��<�j��w�m6�uN�~�"���+���(�+�/�y���se2�����N&y�Wg_�ϸ���2	������EȐF8�k�HY�)0�"�P�~��&�P_B;�T�沈H����zE�7�L�э��=Yٔ�U�<����=��O;�H����Lq�;�e�:l��?���n;���Ӄ�c���Uî2��j�N�_�uP�Q�yy+.��������~{��[��VU�(w���".k�N�����ɭ=ܼ����4˂�f��uk��du����� 'v��K��1�5�Y�>=8ru���
�Q���Ԋ(�wA���!�e��]���G;�N#�iT?��l���1��I�od@h,r�������	?��^��֝���c)A���w��!wh�Ӫ�qQѴK��n������I���Kf� ��fg��q���\9;ȭ2��<���}m~������	;����c�_��Y�!ܖqU+;McV$ㄯg����h�J���CT�Ȧ���?�O�%9T�9�Ľ�I�)Ϻ�4iF���
�9�MGɩ�֝:�kٛ��?��g|��c{�߆�KU!��h����!29�_���#&:8�Uqy�<g}'M���2|�)�if��J�[	�����]�ַY-Q1dZz���^���f�s�[wΜ��˃�W@$t�ꟊ�������+��jk�^�p,,D����J�9љ����v�t���#j��A��~�F��)����J�S��bI��E~�Qf
�/�ܺv�ߐ�n�U�����n�w#��'�%T���e�E�tj�n#mMM��,�~h�?
ixd�s`\Ԉ:ok�9�tZ� �?�oAu���Q���+��
A4�$�	��NG>&���)��"u��"�}S���?����$X6�����g��^_
ܺc
��!TR&IwO��#^�J1����w�6�Θ�x�IG�䒵k��D�y��F{��w�S��7����&���|�u3���٬Wzx&�z�_�{I�IuKD
�g��-�'bh���0*@��^M�@ƴU��~^�FAa�ǰ�N�v���_��gK������S0t�@x���;���M
Om�"�2��9D�Wlpq��Iq�((W,,��{f�M&uƩ���-�����.�%��{+/���ggT�e��7�A�Wd/�ҟ�52���x��
r�쩖�!������>����S ����Ԑ��@Q-~z��g z��+M��q&su!��*u�$������6�0�sz�-�,Lt���M��\�X����#dvA��\�=ͨURw[j�����0�7�Ԋ�г.0I0G��aW����ƕ��c�v�G!��`��Ϧ������ �‛��9�.{��F��K�L��P��� c���R
{x����iT�"9�_o�'d>d�E �:Y�rE"�ʸ%��ɞ�8h��G3��t&�*i��4�,ֿ���]�I�Z�y���������N7�[��u7�Y+�v���v]e�xa幝bI����%�%�	��;�%U�MZN�<W�4rv��2+o�"^E�'m��X�$0Q��@-�U�X�Z�����qV}�95�d�O,��%��Ҷ��@���p�$V�Nga�@UXftog[�)��,m��؂]��Gt�kN��c�.Jk;�Pie�k��X��"S�Ji�B����|T�Ӎ�9�,�t3�g���D�j�U�����(ݞ1,v/�L��i��y�r��r� ���y�� �K�Z����h��Ŗ��w6�gA�i[�]gf����*�AkM4M ��W���4���ce���^&���z�y)��.�����n��Z�9xOy��	h�l�<8v�8<��Lg�5��\�KGy(�_ܳLD��f��:��������W�#�D�KYZsE��%	���J;��E�@/�~Eb[�*��I�����!٧��L�)�#�@i�t,M4Zfv�����S0���ڊT�����ӧ�J���M&ş�ሾ"��`�`�נ*�|��hp�J|F����U:ꉒ�ؐB��sM�^��K#?��r�Cu�Ǘ��G��5��p�$���op7A�����
�͋r�%m@�%O�<���j���pn3���?�c@PB��>�H�߂NN�]+Ȣ#d��Ţw�\�IE�.�&�����8Ə�gϹ�,����d�/�%x�brEt��&����-���I~�U~��1��#��i��d�^'�6�3D̈�s��w�۶��v��/�%<��N`:��R�b�;p�{2��w�RD8�lk'QO���,�Ka�,�?�j�s�fFD�:�Ɉ��ҲY:�(;���v�y�o��1r+�z�8��	b<���x�ͽ�B�,dnmE�� 
�M"l�ɥ�}�qԳ���t���$S�T��U����p����΄i�O�r��+�7#Lm�{>�6�Bo���s3%!�d��Cw���^pJ���J�\a�mp�9�^�9@��ح�z�Ǥ,��5La�}�$|)6�)��;�&�,�ߌ:7��t#x��������э�K�~/8�ȭo�I�wN~�=�Co`�B�	^�G(����s%� p�;Mq��@��#(e-i4�8��
2&O�f$��k����u�dECl0���
��q��JF�2���\kU3\'�,�nE=w��j����rL��g'i�����ݧ����_�I��l p�Ǹ�po�T��h0J���nG����%�ȫ�jN��k� ������76ے.��֍QW4�$MՃ·����qf<�q�n�P�W_�!�3'�'*�n5lp�#�e�N������Z�0�j��$WgFD�1x=�~kѾ����еy��y^��Ӏ��t�ӳ,�;{a�c<y����@
C�]��*X��=���?�mP��R�����x��h"����еy�3��O�U��V�����x�н� D�vR����{�/�n�}��������'�]�ɪf⺉�X<RY��y�1��6�D��T����4H���P��jbM���e��.:é�s�P`/)�>*P��Ga'(4����C����ɨP��I�uͰ�Φ��%V"�¶�.�@km~虲�:7��������1:
9?")�Sօ����՞��|އ+�rWP�:������8Iؓ�e�fnx�>-�*���o�\���ãD�9�:��{��$O�<K��؀�O�P�0�Gܬ���Q�l���>��L_�%�p�7��9��ސ��ʠ��x鈻��X0_1pL������K�i��8�a��m������m�jR���?��g@k��&x���(a��.�I��}�v8:�l��2��>�!6�k�/B�޼�%��hX��Ia��tf�0IFW�����GiGG0���5;���ՙ��
��Am{	� ~�趷u�J5J=HM��:��zbc����l��1ٕ�@m�@_0���.��)�2c��u7xщ��O�-ӇK�5����;e��K�A�[�l����=vP�e��2��Y�{����V8�a�Au�U*U�^�!�RIT���t C�o�<����5dK�]v����0��hڲ��'�!�i��u���y�{4�������[��0cV�?c�HA���O�<΃'�V��wof�Ā���`��+�SA\�~�~R����Xi9�D�c$�k@,� ����T������a����=�9���M���%� �U�̳R�[��ǃ�D�1ڇ�1&�4�q��6�ٞJN����),��	���5�����iU���Y��k։��|o�6ѻ���X~1�@�q�-�y�K�،����\&�������ɦ�b�s�`�2�얰��hk�{1� b&�g����ө�'��؎/�ܾ�����{ĐD�Qp49-�-g��^M�����b��:�ml]|a�d��<�ʤ��"����ھ�-.�^0���=��?�Q��TXطnv�d����<�➀�(�Fod^��y��ԯ�z����{I���3�6��=B��Y�ZQ��6mxk�Vm�J�c�wL��k� {.I�U��y>��P4'b�dIFl�n���t��z&�C�X�����o�����r�/�_�v��D�edy��_
�X�d3�J�f�=���.�]Ӽ*��YBam��s�,;�)�Z1�!���������ꎎj�R᥃�tE�H�����1b�s5���3[8)�*Hw%��!n�K����(�}�~�( �c��s,p���m����L����&��h$8%�s�&z�o�����أ�=	l_tݭF,�jfU*~��g�#��_��'�$�ȶ
>[x̕L��e����E�u��XG��ʱ�y,��Bj��.�~㨷/6�m �w�ieŖ"g����J����;��%`�� ���9��%ײ�"����Jn#��o&��1yO�q�Cv��0ҽO|�ĩF����nBP��,|LX����⶞��7o���j-�7h2H��� �1Q�S!�"?�Tժ�3 ��C��r*;#َ�?�2,�[�#/����1���o=��%PY�hʸAR���rv2�p<�xd��1�w_��x#p�~�kk��W�)̫,��&e;|���4"G���u���^�lc�������4���Lҁ�~*^��4є��Nyh������q�����&p�Y3��P}zH��	|yD�2���b��]���m�K�K���>�0������6��r�W
�o�c�Erh�ɭB�Z̬�Y�������'\�۟U��c���%֩@Xo&!�f�d]K5E�::=�H��d�\�36��R-����2^��s�J���U�$�W���9��x�O˭�����]� ]Qo��>�{�r%���h������������4N��rEJ]5>ѫ�)����O'yM���|M��\����'���6ya"&r����q�pАG�3zilhbt�+�99^oȔ�u0�HOά���(R�G�)(�!�c��>gM�q=r]��5���2�)o�7[����3��K�Ơ-�ƅ�IzݞU������V��"[TH0x�:g�㿹��i�a�~D����t?��Ә��L�`7 !>�NER�K"r�����u��~^K�9c��VA�5����M]�DO�̳�*��A9D6���;�N��L�G��}{���P��u��	��J��ڿ�_�Ѳ��[�[S~�9����c��V�Sr2�p��ŪC'�h�^7��h�u�c9G�����jtr��tauOɖ9�!�y#��U��#�$�W�ePH��=F�Hu�R(/�S>xd��oɶ�Z��G5�TA��l�bi���`��y%,Fi`�� M� ��>��E��y��*s�*o~J��lI�J���3+�4o,G��ku���.�rS�2���b.Ӗ}�<�S!l��9�/���H�S�&�`��P:#y�z2O}�X��#y�dc-�$ʒ=�!���ڪ�XR�Y{rS�� �˗���(aJ �#�>��G�]���<����Sw�ϙ�da�����X�=EX�t�����8�O�h.�t�����^��� �=�ҝ�)iBn��wls�@���w�E���^� Qq�b���U�|�6���c �u#�&��w��X����:�7��]�;Q�l���w�HMgVݷ��٘����Oj T>ѕ������,nm��s̄��.=W����We��� V�C�ީ)��<e<�YF`�U�����z��5�v�u�g��L��B���^�o9��$��n��IC�?#7����JH��rh*Z?��=���Q��}��0(�]l`�h��Z��<��)06����C��1�67+J��4y�{���L��M�����2=l�b��є�_Y�}b�eyK���[�	g7���i��iP!�sf�wO�o�Y�K���^5��Z*?ϾF�#H ������r�ӝg�Ql�wI�����^'9GQ�����m�;b�!��߂?���o
��<�ߦ!2�=���a҃�R��wZo�@v��^�����=aT���UV9H�a��a�o�Q���y>%L��j�{�<k�����c/�bv��2�Q��O�ؓ���,>c2���,�[p��(�ۣ8�ܪ�����ܳ�8!'� ib���)����/�9c�ź�Ⰴll�8H�Ybԥ7���Y���)��D�n����ewpR���3�#W�ǡ$p6�eK�Q�:UX����Y#��#<@t�4���g�.�D�n@v���f��G�]u���D���"��Df��f� ����O����$/��e�oV�9>�R�#��Ε�i��?��>�Fg�-�z�?�kE��o�a�"�,�(�`�N�O-N�9�'w��n���Wx3Z��ˉ�S�_z��3'�;&N	���Uk��a'�8�������}z\�}��҅�)9G�w=1�@�pm�����������j� sP+ĞI�{�2�u4���d�����%��Ί���V�R���������n�6.Fm	U�7{@���fj�x���G��8\c�,�Q �$]Kj��/�������:8_�0̲���&�iߖ���O�#n�d�.�uCm��n�n��s�$=��
?j�s�޷������ZbU'iI� ��ԁn?
Rp'�~1�.�T231u�k�g�ި۹r��kq���Bѽ��aĻ����*��4�I8�@L�]=��h;q��3y�4�kT��Z'H6���V0}�ѮWM��7˘1פ�V��G��:怈��)�q0�iKŕ7V��u��@�.�n�e�@笄O]�8ox�Uԥ��_���F:����Q���M����Gj�u�?7��v���u]��Ur/��o�=wy�Y5���ش�9�@��#�;^ԡ%d2�̞�8׷/a0��㣧:���2z���y�|�o�	F���tj慨��N�2	J���m�_>���.)V}��Ţ�x�4|{�����{s�d�K�ƶ��woLO��2�,A��Z�9���޲<7u���5:t���X#.�&��x�1 vFI*�6G5*�s��uT{��n�%tC�Ң�V("BNb��:C��5�<���gb��#�zĹ���I�ކ���� T$���x5'�R�Ms��92����q�H�O���������lO�E���s.���z�h���r��
T�L�����%���O|Lb���A��7�'R��k�Ag��p:;���4OhR���SS;�z�����"���X]�^�i;���SkgyIR{�'���,ޡS���4=��zu�s2e��9�U���#����\\�<K�����u�Sl�2�i:d�^�M���xgKЍ��r��İ��P;�T9�v01�ot�%�>q�gv�c��4�b�\��M�R�<ƅ���(���#��Tq�{G�5�e��� ��h���W#�������B��n��R�,��G"���1r0ț;�w�A�����;���3���ܕ���e'3\��h�a��;��2�!9��_����S,'!h��*ڞ=�����׭��'"�G;`�����JJ{��I�ᓙu6.�������x!��,:T���$#l�w�4ZKao�vBq�G���|��Q���,�#�=Բ.\d�!������u�R#��c�t�T�o�[�@���n1�q�Y\�-/��T�(��{��>1ڄ�',�f=%}����ǹR��%S/�/�$�A�{�r&jj:���������h�z�=h�aY���C��z�A����А�h�76Z;���	�s^7��@�.��e,;Ң L����h��N晉��}Έ%��?��/�t�S�]�Ǝ��ͥQ��𡶡�<\�V�E�CR��~UkL���K��?1M�-�ɷ� �M-I*��I���L��܍}�n�QTy�oH�=��Ӫ���T�UW��a���d�oTR=���1R�Or-U�}���ĭ8n:~j�Su/V����H�"�T< ����OW_�J�a�
��e=R:��5�p��[�,rɦn�Kς��^!��n�5w���7����� j��xcml�����ve
:�1�;!�����J��Y����n�
&��%�y0~�8���1+� 8��.I�+zo�/57O훑U//��H\�#��G߁�8Q����^|+�[Msi���}���ӯ5@{w�]��S�c�p�N��d��ʈ/ÔHA?�4��O텴�G�u#���V�e(��@�t[�\8�X8��7	���[j(y�Oմ4�9Q�D)Uf�I8���w~h��TZٜ��*�N�8,?x�/!@�ù�[����5��t�t�j��~�Ī���?�w?�ٟ2حz#�`#��H��Ov.��73�7��@��RU��pC{���*�E���q*�cl�\��V�>
z�q(�?��������P�*)�������=:�K�5�'P��(�F�RO>���ޣ�:q���ϩR��o�R�sR�4k�Aq�`��w�v<Yp���2���p��i�lYúp�.˂��I�.6f���ʗ�L�gG�ֳN�id�I?��u��5��Ag��Z kW�^0\�%:�B?�Ti2ruӮ�ɑ�M�PM�}��i��~�K�<g�Ī��<@�5�D�\'d9���5��X#��)A|�}H��9w��N�z|�.�2�,
�(��9�M�;W$�q�IϽ��8��'Ι ��`s#3��t�ݝ��EU��<zz�Rlh��UXI*�7:�ZjPuS��rp�Ɩ?r.[�K����@C�u0wg��<7�"�w��Z�!t�+L`UzG`&�׼�N�C��7�|�=@W����������%�`���.�Z�����������S�Ӹ�.B[�t31?��r��1u�|��Vu��m�p3?�m�e��5�(�����j����l�*��v��	:^�S�<P�q���=&2z^������X�Vt��<�Jy\�3Y��Uzm�㕒1�z�{���݈<���T	颓^�^ ���Z��1���4�ᗜ�}�װ%E��=J����<��r_��[(g
U���,���u����$�P��y3��X���U-.m�5v
=<�OR������ڻ[@:�a��.���o\8���1���ץ�!p#ƛ ]R���m�)wZPh
*(�O�e����lh��Wz">���X!��S(�9�57/
[��}I�MHʕ��|J�E�)�x�	��B��'�T��Y��Sq�s�KMYyNA| �s�dt�a�G{��Xd���PՖs܈��Ҥn�aG*�a��7�{Q�r�.W"�%S����GO@�0�"	��=��D����O���}�*����ҳ��K��o=�Q��)
�~u��9b�>����<��qv���h}�q�e�6d�52-��	���"싽��͕a��Ǟ;��NcLPz<	d��G:�=wt�|�<�{���
����LR�l��ɍ�U��L�}�Z�_��'��vR�&���j���L�n�yU�Ⓗ��Vn]l�;��-��[g ��&�5R7��j��0�����)1>�/�*�zoE�8J��������|#����p�����c��|��JV��[zc���~v]~��U���ڮ�.����cM�xՉ�˾ʈ�`�E��
�?(s9�	ֳ�ە����}��k�ح]�� 3N� � ���p�?hpN�we������x@��{ 4τ9��-x%>�J�$ �-F��(.*HN���f���#���4\�&	�m).B�l����s�"�Π]�5�N�!\e�*lhʝ���x�<� �|�C cY\�ńP<�䨒���NF
�Q�q�v��mBk���m�o�Er���P�T�A����G��1�҉a�+`�6�(�$�G��s0e�],���P`wr�ϣ`�$~��2H{c *xĢ\�#G����ZoH�H�LM����IqW��,�<ں�ۉ}f�owUӊ;�/&����Ş�#������l�%�SR>N�]�H�NL�\2�܌���xC��4�uŇF?��\5Cs*��H�6�mA��FL"˽������|���!�!:�K� []�� ��9b��
���
�l��𞐶�VQ���]c��רz�q*5��gg��Z�9��d��x�l;k*������l�jo��E��5��@8ύ����bu�v��y u���(�r��M���7zƞNC�80Y�c��>Q��~�LѠ�;N�`�u�6�d�H20�]{��q��^���ԡ�b"�{|���f]r��l�/5�,�is��h��;�K�V��_���<;TĤ�c�4&^��K�O�d�Ҕ�}��-�E������"Q墟*��}j~ƾ	K�����c���F
S�>���cV$�Y�ᖮ�ZN_�ݖp%���dv�տ
d:}i��nL5_�Sjԓ(ڬq�W$�k*�Ӏ���3ht�����=�G������E������v�XC�H�N����I�^�_�<�9�g��>������Ȅ����@<�\�9g��'�1�4�=������.~쯫{#�,��0i<m�L�~�2��@���:��3�MPO��7R��ֽy���.���|6Z���_���: �ݵ쓘J�uϋ��>��@�L�y��lk�ZW�gb���\�J쫛݁(�稞������5��S&�yNa^q�s�
q~m��z�/�\�z�p��n�Ǳ_L�����4M��vR"���6��eqa4Q�Ӕ��^V+}��>�ĵn��F��碉߃�WX���Ğ/Tb���1-�����-n��4�V����X�L�F����8@�����1O��!?�0?���
\���?6�O!��ݙ��ķb�A5_�kB���
j�g����i?��� ���w�\)u�5 *�;å�R�ַ��I;(1H���%/��v�V��D�CGl�c�`X���P}$�\$d�D�?����l���^-�Z��5;���h��den���[��0	�6�� 
�x�/��O<r�v��,P&�5m�p�g��\G^ �ĭ���y���+#�@_�Sow(5�Q�Ң�����@�$Ԯ�� ���\�jV� 0o�u�2�J�)�a�o��X���oJb9nz�z���]�e�F黾(� ���M����~�.+�����o̤�3y-I��Q�m��>k�}n
�'&�$��h|�a�l�!�B ��ܕ��yUV�]����G�î�JH�jd�Q��kQ�_�w�Dg���,xn��Z�7�(g�
�Ǯ��t���3��������!���p���N)3�#V����-T�OT���Vo��j%�Y<���i���v��Mflv��h��WKj���a�����%m�e�mP��G��R�y�x���I���n��eu]�����ԯ��M��i�D����~��/9Q(��2ほ���t�u$�P�u���)5��%F>r:+��7w���y����ٺ�;Z�s�LĆ� �vNm�6T�1��e��3߈�g�R�^�c�{]��h�n>'�x��L�*m�~c�N8��u�5�}�,�L;4���z�DdCm���Sn�b152ᮍ����'P۠o���`�����=A��z�ϱ�u�_��[���Tk���3�Y�ꂴu�s�����P&"nca(H���z:��a��O�^�ji�M��i�͕��ZQ��a>h��6��C�,�m���i/��%��#��8��I�D��fW��s��|A��N�U2k GW�mT��^�e��V��f&t/d���0o���� ���+m��該|��!ef`_M{�L���_/ʕ����ޒ73�٪@���}�y��Hq��NOZ�U�p�s.���E|�Ppo;��� Y�S)��Q��r��9�N�S���5�C���fpd��+#�N��0lႥ��Ģ�P���_�)ȡ���{H��=c�#J���#ɂi�3�;���̠�!*��N_�H��f_S`�v���;%���:𡔀��8�\>�*n7��%q�171��v(��u2ԉ��a/.�}3��x���n;T�ql*Q�F���.&��8����{
��1��c�'~��?=8�W5Bj���{y���|��3���/�<����n}2�uЁ��S�c�2�3(()����K_����ܣw�$�p��s�.{��!��"�G5�W`h�܏�Co%�v�hKSr#��8�:m/�u�"�[�[e�x�Q)[ddj���WG�q�$ɴ���뗰�Q���XmZ�W!��8f��[bb|��x��i��CN��ߕW����'髱���3�:�r�� �����f��c�-^����*
��z�)���e?k
�tǪό]:B]�\�(b���f���C=c ��b��0�LUNI���!n�d��%]&ܷL�Rn�;ɆfI�I�,�l҃+�O�đ8�f�!�>��&d�;�^0h2׾�.��R@I5K���w���y��t��ikY0�B�L��v���$��g�W��y ſC�3��"�B���Pd���Rh�_��6밤3�H�Y�q5'O
��e���r�~2���@������0�T�L�k�UqO���mVLPЎdo���M(J��Y���1(b��9�pWj
)��� ��<����}�Y��7���$^��b� �pu]�Q�n1��[L��0���рO��+�7��������u�G��M�*�i5W	�M�VlJ(��vb%�z�ؓ�����k��$>MPL�&�
����)��w���c�^49N��7�I
j��L��8�	�;ܒ��I7J�Z@��_����(��RR ��!�}�\��?�g]!���PE K���̾a�!/�!�YD�i2� ������NER����k�Lm��'L���I���0^1uo�Cn��pĥ��!@����$qG�g��VL9�c�ji�]�qV&2uMJ1c��p�O��]ʑ�� �\~�F�=,Z�[h�׭.<��B��a�\X�֝�5����LSb�t�,�M��s�\4�����C�6m�5�s��D(wZG��Ѧ��xF�� ��B�
�sv���*HW(
'��rP�EZ|������g�E$�7n��������t���`%���:�8u\l���t�@I�KF^� Mv�CmNg�<���]���s���6E���Bv�x[�[U�����̳�G
J��p0�|��`�F7mv����1Wq���y掲w�9Y���QЏ���Td�r�&gp6��� 0",��ӨaQ�����;O�jn�7Ȣ#�6����dnީ3c7KU���B:'䑡�R�i�;��ձE�f�UaZTK��v�G�y}Q�Sj%�4L������y֎����=�U�JH.zL�PO��*�ﱮ�=��q�eZ^��/'����֖�\%VS{�=�	9��]�Q������d���8�YSiMBK�-��M��f`�d�͋���DAO~mef�k�^�2Y �������}9�U2�!�R%��+����v���a^�f�ǻ%LW5�=l�sP���M�����K)zJ�l,,�5�c�7HS�91`��1+�Gȥb�ll��D�V�GZ�l����jO(x�&�Zj\Z��/!����R�,T�x�A�,Yp�����P��$%m�͏y������G�-\?G�FJU�GU
7��`�]��ΓR���)d�H�@��CG,E�Q8�RF�9���6�Cr���ÎRr�δsy.�����Mΰ#ld��������)N�*��O&m��x�<U��f��z��������a���)�M^��k;�l��2����bFy��8RE����2���v��#�ˣq-��/>St�z�yn�"�U�L��R y3R	�Y6��$�
'�w���3���N��x_�� ��F���]0H��])��c �6��
��WAol� �<&{�"�Gs�|xm��Q���ϯe��uQ���=��AB���N�Yw�-�_��2LQ�={���x����Z��R	w���(��4H�8W��j2 ]��!rN����(��Bc���� y��;46Bs.��!�d�e筷q^��6n��qf:����=M�(�n�R#9a� jN���&����*2k�l��S�'���� �mp2v⿜��|�d�,���ݧݭD��-մ(�|p��!���f�(����^:ί����hS��6�w����1��u榠�ڢ$��	���u����O�iI[r���1(*$�>ҹҞ"�����h�����)0�%�\���/��b�Qt�1�aU�G�	��%�u��9���!0�k:�F�<�{�:֤R�L�~.uԠg�ְdg�
�����|׷��=0�X/�pT��SB,D����;�t��5�f�l�܂�����;Yb�YV���u��bXP\t
ķԕ��3n���O��̢j������[��a�N���!u"�H	�=kS،����%OfbO��)YTV�Os�lY6��g�>�K�Ȁ� N^�"����b��C��4�b
"w�5�#����_��b���'̡��o���&)��,r���#�T��������i\����^VHZ�Ȯ�%��ڟ+J�	*\���rW����HwcG�WU��S�n�qv�5�V�U�����aP`�C�{&07�i�����U�}2*��P͹� 1��?�Z���;��EJͨ����f<W6���&��{�;m>uJ�&ҥ�Φ�%X���&����.�#��������!ED�^pgk���O҄�mގ�\�w��<-i*RX�e=�I�	��	w�Ҏ���}X�,�QX�v.��]��S�e�}�Cn���3�8�!l���DPc�[Л9��(��A,���Rfv�j��<�[-s(e#nJ���4�� ��'@\�7	:c�]³_wqY]y�W qC,&X�P �^S���)�oʐej��������겡%�G�¸~���c��=�@��s��t�{ђ���=����P2�����̉�v��)��H\0�o� k��u����0V�����c�/˚�q�<��۩��B:�D3���Pǆe��ڋ#�09�'��Dc�v+�e��N�1Yz�T,�l��%�zI����C;=U~�i�u�]��~���|%
e *?���6
�6���b�\�M���(C�T�^}P��A�N��IQP�LFS)�E"�l�{��^�iy,���r����/����;���n��CU^��r�6E�w�az��,WC~��m�:�Ų�֏U�q��,-�	/(���x@��p�����`V��H��еy��bX\*�y������jwY^^���Z08a�mi�@N���k�؃x�e@NW�)n4W�v���BX�F����=�%v�B��&ٱ�� �jw� Q���Ms�+�Ђ/w��p8����;��ak��gq������/��@8-��m��34�}v���o4���v.��V��N��IB+�r�Wk/��Z�u�p�F��9nu�dgڿ/F?�Ot�d��-��)���z���(�|�HhM�A<�{�؃�����e0�׉J�ZEg��)6dIG�}��0Ynz�P�Vw����o�ڋL9��L�f������60|� :)�����Ǜ��+�^3*s�'�*/��$B<DbP��	�m��(%��S2}�����e2�]{��9~�BIX�v�ZS��g&��5\_`�9�����"�J8�"j�QY4��Hf�p�s���t����#.x�A���w��[�I����g�4uh]����7�`c{�d��1/)�� �<�Ŵ��@�VՈ�j��EMAya\䂑sO\�CǇ�	9eG&*�"��ӂ����SJ�Vt6�"�/�IK����K7�?�2�JW3Dܝ�^g�ݫ����wGE0�d���]��aZ��g��A��j�1��i͵F�U6��!�����Xʡ��y\'I<�A�_s��y�-0\v��0���F����]������BJX���t��(��u�lh�O��I��A��Qɰb02/5|�Q_������h)CL��@���{d������M�EZ�g6�hx6��R����U�S� /��Z)���ꌂӬ�n��w�y���Brn�	Y왣g�l�>����f#�*�Y�%;��5���i���!	�{UƲ���rr.� =�H�66vO���ΏW]�r��M���V���)�'�8����O���WV��x�0�����	hy�r��&gP|öt.ܬ�dpߕiw�O3u}��Wݵzg5���NR[�;�����rx�����4
�L��m�<d�*��T�Ǔ"}�[%9���Yl]���w���Y1��W�%��n*�t�y_	{�6�߷������B�aS.���d�i)�Vy�eV<��l�4}9�|�^̩zr�©�t�zX���ð���	{w�[�*J�{K�>T��Л=�1}�]��KZ<B�jP�'�����j���ת?��;��i_]�ڈ����g�K�(�tkӒ�q1o�Қ�7����3R�y�|�^9�
S��j\U�4,�$�7��Iro�|y2|&�����2��L�+��5[X��~j(7A�A�6�Ǎ,����P[�<�����5<S�o��L1a]OiD��x�c��r��ܹ���(���$�8���#��}�f����nR������8�|nDW��b�oE�+�G�A�Niz���D�z�r��H�2QĵRB7����������_�NoB�CX�����u�Q�����FiA��X�XK�H�:0��r�_�'�%�
�.���i�C�(��M��C�]Q���"�n���P&]���Mp8��"��qwt��i+�d@J�o�*��*h@?}�`�@D�
��W[+e��nf�S��pt"��`)�5�`>'���ݬ��R������T�Y��_�3�����^|��6�Um�߰�>��g-�QI�8�?�1:}$�f����7�%������c��6+S$A�1a��D˱k\�d]��a��*)���� �ݠn�W�(����i���ð8�M#&����3u��(L�E������h�㇝.W�/޼J� �l?V�=�p��Ёk�'}��y�_3��s�on���a+9'o�g��o-�D�����(�|��[!=��F��V�Ka9'��񖬃ך��O��H�A*�'��FT����a}Aa=��ϵ�_qwcH�!����u��p��<��X�ӳr�)!�9�'�Aպ��m�?}s�`�>��v�>X@�|�d0e�$O��y�cj���>�2��d^�P��k<g��շ5�>��a���T�Eu�!�]x|�����S�Ks���*,]3�BM �����jx���=�"��Iֱ�%� �-�թ��̯8Z1��XL�#��rwO�@8��#$8�Q-sJR����:�y�r���(���'Tz�xDwܴN5E}{�.H:���&��q�c���ba��>L'�4CG+��K�3v�
�Nߜf�~�q��j���o�Wg�)�9
qu�����w�|U���Lp��R��^+N�n�!li�ܙ.^�v�*ܻF�$w#����,y�a�N��s���ª��4_;qҪ��غ� �g@d�$Wڧ,�$Ph�6;��mn��?`�sW�����%���-�����{���z�mm��d��D���+����"CRCp1�����8U=X���VR!PR `S�b8��l�?Z*���W�(�/���c�����H��O�"=��g���o�z���#⣨�L��p
<j��X�H[p�Z'��Csm��Ӟ��gN��-�N)��~D�{�9#���Fy��2DN��ѦI���)�5�[�ӧ= Qee���I�;�R�ٍp�M�n&r���-'d�pN�'���gG)�8T&�P�U��<��2�u�O$�H���W�_���f}��Ϗ�^�jj	�Ԏ��q���*8q���$5%ʥRPM�.ӼN6(r�t��.7�����}��%[��uQep@BJJT9dݚ9j��Ʒ��ʏ�ܸ~Ve,*�P	[�X��0���ʒa��W�ˉpx����y�r�S�. $u0R�]�	�*�S��_�W'�6��Ċ���v?`�C�+������K�C��ޱ� �'wE��}��Q��E(A0�-*4\����n�A�ަp���ȵf]�#��ð0hD��.�a����Ĝ���U��ߋ"��c�^�}��b��rk�
'8 �
b;�h1PSޗ�/U{qfM�r\��^|���QbC�K��B�7kQ������ь���<����p�?w�Y�E�R�e��Cz��?������_��!MC+ɾ�a��,�q֒���+:JR�*e�k�FW�_���GOg�՚���s岚������:���ˀ�λܳԤ�a�oE..C��O��@�E7e�~���+���4{���&��M���ʃ���^XE�\�=�U	�P�hv���"�>?C�����ݥ����Dvw��G&,�-���!���qȽ1�v�tAG;�����[xDm|�O��v�?OV鲢f��A5��/�fqO	{v���lB�M�ʥ>pX�{�Bu*Yn��Yp��	.�hFf"�3z��{f�V!�w:�ѷ�}����JֻJHΙ�?ۋL��o]{%8ЍD3Y�W%]<���C��%�-�%U�欥fuM��ձ�Tm�?�D��X���J©3'���~�f�Wx��FWځ�i(���0��'q�7-p[<X�����i	��q��N����C��[BSN_	C����}%!8�p���
�:��[�V�3���>�P@�f�Pd��r<��8m{��N�bj����;��b��qz�QA���>�␉(�1�)3NnP^e2�)K��3o��0�4T��O�5���B/�\��|I��͚�b8b��7�oZmg��D�d���v�T���]`����!&��r�.��9*��P�a�+�!*Q�ɍ]\�w{�x@ ��U�Ǖ�'1V����Pl�y+����-��O���u�9g��͠����E���x$�~CK�`�>#qO���a�k�r��e�b �І���x�Y����Cl�K��3��l��`
K�#GhkĮɮ����6(��;P�\�|wF����u��J�^W$���	����1=����ĝǰ����nu�+�r\��+\�g.�j^�vh��_�O�y�p�9@�;�J���i&|R�DQ�ki��7�_���+wz4�o�7��H�g�%/����sք�m�)B����K�0z�v�(�ά��e���8����tR�<���5���E,�p���qpv"ס#�u����}c��ǆ��*�Ĕ��J��F���/��u�-:��S]���'��yX�̓���,H@��^gF�b+(N v�v�<�(4;#�����íz��ܸ�q��ɇA n��)����Ǩ�w��;� y�>�>�z�C��N����Z��}��B)����T�� Ax.ವW����8h*Q�{�>�U<kB"�|�ʾ^����կV-�����û�%h��9���cz�ai'�0yM� �g���E9KP��٤ q�o��NekJG��8��j����jd��@f�G$O1��L�ט_�,��
��Pq�:z�0V}O��Hx;��z3&+�t�c8� �s ���o|v�J�$R�ѥqDd*�	�vOh:|�-+�g�a,x�����ՠ��%sG��9�Gpw~$.&>:W���ˇoz|]��r�K
��Φ��w�=���$�Վѹ+��b��U@�	)!l�c��1���K���dD�O?��t�+�.�/��mJ4��u��%�'��.p�ؙ{(� YA��R�%�|�|d��Y[�#�����-�j����R��$O�fx�}�i����-�ߴ��<	�	Ӧ�r��=��X�%��PC��z�s�v���r̉�j��c����VQ��$��m3�bPVI@2w����Oƣ��t�}�T�f��nk~���[���ɧ�М�R����=vd���g��\����o�IK٪��3����(b�G���K����9bZ��6�7u:�YP�����*tH8�FJ����R�-��_�"eU�K��T5���WI���3@���oT&o�'��˥�&>RH�od1ͥͰ���Ct�t�q���}Q����V�G&��L$�����fT�<[��)�T!����U�7<�"za	��Bmy���0�?�8�U�擡�Uu����C�w�6�[
�'���uD}{�Os>�1�t�ag���\��������D�RkYe��L	�VU��	�È��+L����yƪI���NQ�增�t�,�H��؟�q"����PGH>{��H�� ��]�F�"XD,cX�|ٜL���I�.1����ƕ�l�ޭegS�ػ9�/T�J�mEK$��R�����W���� ]V�*g'SP�'���=�%��X�Ǟ��nS��ͩ�$Ih�-Yts�I�ݝ7�'�`�*6�4	� ����8iT��aAz�gA-J:�c�:�
�F$W�� �郦�4��̘6+ t���&�D�l�jƵ/�:���z��Z��M���C���������	p���goQNVJKzg�5�<Ef��9^ą��εX'�'�g�C 7V��R%���5N�~�J�e;~�r��6��
�TM�����y������:�g�b�E�w#���T�I0���[�G�$�`.e@Og��*�|�<����E"&�~F%��8JI���/��\�J�/7�Q�~��MmGfR~��)(�)�S3�K�U�ғ{�c�<C�֔����X��-J�\�w�z]l^�H�3���[�9'���,�_�OT�e;�ӯ=�|��]�� H�-��oCX'��O����H��^���f���Q&�w����-үa�!��,�5���/�����ܗ-��� �(OZ��$���a�(�����bT�PޥKŰD���N<8�:��K�PvO_�T4>���FR�DCG�<��B�ɫ��B�O�����Z /V��������_+ C(���烎��v�2@��~�������K��qf���|��h��=���ѫ����t<��X:��S��뾏2y��K����<�i}V��1[MX���qU��J�����A3׈E�Al�W��ۘ��9S� ���/㛲,�*�šNw9K��D���T���H�Ɠ�F�>��t}��9N��1%�uw_���`n_����MR���q�i���P	d�>�.K��� Δ�:��1�y���t�A���r�?��ho��
�����_��\_���0ܓ��n�%��~EI4�h,��%CѴ��N�<Ҕd��oF��wk;��$��t��M�o�0�u*X�qF���E���Y4H�M�g#u��r4g�8�Udz��HR�88uV�S��6d6!��;�ca=s
�������-H�������۪o��!�]�濞a&�jX:.���m:	BWm�����EK���F�E]��@�����$�9������ �~�����x`���;��|U��8��0���T-b�j����z�U3fudpQ��mdCb���9Mɓ�.2�C�|'�@�=������������g�v��i���<��5mH��MY�M_����4$����a]D��(jK�R���5�vr�4�(l�u�?#�*��%��M̆�Xep���C�1�G2"��������ە��9h�c!�>����I�ƧƗ�B��X�D|h�#�PLdM,�_�&��)1�Y�����iܼ���j>U��ܪXmȬ2	o�H�b}?��Mw߮,H���l��2u�_h�pL�س�Q��7a)N&����a���yS�}�"�k����Ǯ�0i�P�;����D�-�P�m_q!�W
�c����Q�6���C�9�W��C��\�>����]�įߥ�g��}��7�t��+��l��/X�˗_�>Q5�/4��������ciI��[m7��8�/(t�f������Ma(����{~�MQf�7=�;����U؅�#����mH�Ne ����|݌�ƾ�C�ƺ�=x�6���I̭�x�-����v�i�^��{ԧ>r�Q��r1Z�=��;������UVZ�<Rh�rn�M�ߋ@�h3�������16W��<�!���T֛]?�4'T16�H>���[�5�6r��[�sm<�s?@[1Ei�=�̏^4@,�� ����c�n���\��3J<p+^p�	O�g�Q�qg��]|0<K�R�wB�U�~�jJ}��E�5�!�j�>�A�0�����������3DU��}s�X@��J��f�uU����H�8~9 ��jZ������a��44��]m�A�ĆKǷ?�׌_�J�F�o<��;-��簨`�!�� �+���W���\�A�T(���y�_}��V�V�M�v���E�f�w��~��4tS-J���Hq��%\W��`�RB�,;o�b{��_cxt���ŜW"A�8E��4H3���"K[�G����u��dQ���Ƣ���bJ�rYJ\q��!��%�dy/��GE-��_��Ϥ��BX����k�<i��lA��[|���Z�.���v��Hߵ`.w��b%uA;!;I�I�u��ǆ��]	,tA�]����[Ĝ M{e큊A�@�{Pv�H�\m�$�j��)@HZJ���s��ψ�>�Kn�"�K�T�c�HSZ�Xx����'Bw#��s�ȼ��C��.�sY�:���5Nݵ/+��m?�
�V���\S1�	u�\r��ouKn4�dRz���1Vni�����ݏ;,̐T��&%)zV��pE��ڊ�nWDh��6�p+�lڢ�bZC��9ւC�p����i�93d�՟?2Z���S��)��V�)���,�ԽU�h�3��܆����~�Q��_�:�|����N��0Gc��7A4n���Ѣ��}/+#�]�'� <�>	�01i���S����V�h����8#^���?)mlX%���\��Z�#�b.��x�L�
�i�����W2�-e6��ĕ}���Y���"�ѡq��4��]��\a1������ǝ_M2��|ҭA��8��;�>�L�.u�eU���}	D��XM&��nPԕ_R�yގNU8ǝo�رG�ʫ=�7$����5��`�0�t�ߧ�]�˩� 	�����Ԅ7�-۲-��*e"~`�WR�9�����2��	0ЇF�������Aҧv/Ԁ�VUe��̢�dv��ʢ�]h���2_���|*�Az%��$������"V�XB>qm5����`�{ǔ��S��Y��u�t?_8��I�we'Q���U��V&��Z^�u�2��A���*�^�� pa������{"_5������<x�1��qv3+���b+�{n�q%���p��g�VZf�jfm>�v�.�;ihI�`5�{k,�=����@MY��8�;����R7&F�k%[�4�@�t���D���d�y�4A\>��F��G�/Q-n�]giϭG�D4pfO�􊇡t��D�<��7]�gj�z�v����Go؟#KdX*���;<nt��J����)��&Ѡ`1�oF-�������/��N�/�u�l}����4^c�9W��>:����@�� �,�d`,�"͠:����ƁpJ�p`�I�$E	����X��,�Mb��Kс}�2�k��;� A�f�6�N���y��@�#ib=�@����#e��r:B9!���Ju��z�����cb^�?���ۑ��F�f��v���%�A7RZ3��8�)nd8����C8����|%Iz3���qͬ.z�
F�猜M�К�t)V�	�W]Y�y���f�P���ۉ��`Yo�k~q�굆l"�\����t��^�/1s�����@�m�~���l�'u��?:<Q��`s=Fi�!�"�ӷi�b���>�r�U����7��v"���WR'>�Ǟos�(x5G�,�jJ3���0Ͻ�X�Y}�`�����N���Q�,6��bfZSj��ȑ�VqR\�Q�jwY��!31�X_Pqqt�Cg�yG��t=/[.*�c&b���D3-_��n����S}��OV��y��H��/8�"W�6?'��M=1G�j�����9�N�c�5d>۝��R�N��&�����t�u�����\e�?����^rK˧$�1*^R'/2���dN��Ns+V�0�SB��Z��n�KL��&���_�Y)�v�����#���\0�`/�b��GsBD�H�,9V6�����Ǎ��3\��������;�ޟ���U����ve2%�\a�Bh�`ݴ%�f�����#q�Nza�;�w����Wdbsn������1��;(��%7������x��X����	D/�Ĺ��`ȚZ���N�k�V�Vj��(���
�"��{Lb��8�ז�ef�����S���}EE�ᶇ�2pRcv�a��%���_e�Бv�ӻ���!p�ڄ1ڔ��nV��pXU�6���,Ik瓏%I���^�3��؎j�ʧ��y�F�Q������R�о��h?a���z1o�f���uތ+Qg�?���Ȯ������/|��Q=��R��z��D�2�ލ}�}�N
t�]����`�|ᐇ���}cERc��"�PT��4g%ư�����te�$0��ì���.fB����|�ml-���9����a�B�&�Hk�(]4Ɖ��n�Y:.ư��hI�*���.�o���p�(�N'�odH9��g�g o��YQn6O��2�p��;쥈��z�8b�G*G��`̿����>g*tK�8��]�(p;^g'3���P���ؓ�l����y"Aᩙ.��f��-�M�$2B�&�|�˚ڃS�����_I�(j+V4c��jZ:�òX��=$�p��{$���&N��3�z��ۼ�ԙ���� �-���fI�F�Hy�ìY�tP�:)jbY�3�!�z�N����z���=�"�iQ����O�������[�W ��JG�`-�wԂ���=%;��QJX_��z�
��������4b���khޟ�g�"��aKt�T��S��-D�bWx�"� Z��b���hCE�!�y�<i�aϼ��[n{�?�椙�@�[��B�e�6~!ƾ�2i����e��]�qNb7�k������ʎf?5:L��u܎�4�yo�W�0xW� _r��q
���R}�_�x����7�1VA��G���t��xL���=y��:g��[�AD���Z�|���m��\��r=.zd����.�-Iǹ�A���	���z�� }+?���f�b�]Ҵ<�f��<������f��n�y���v����19^5�,H��ҭă��Vn(Ԫ���d�R�KXT�j�#(��x�q����K;�v�j���"�{��Ļv���T"a{��JŐz��g�����g�pD���#��0>^��`;��R(,Uh�>D�J�)ʮ�����Vc��	X�d����s#z����0ٺ��t�Y�#�9��m�=�M�b<���	�||H�Y��1��!nԅ�+Ax��k����%Rxkz��@ag�9�@���~�0D�=0�w�o됮4��r�4ƞ�p�@'�����zM(^��z'��eMNޢ�_�ȭ�n83�4���;��`KP�ί���<u]9،���.��$,�6m7�F�#��ۨ�z��G� S�S�}�1�a�Ю2cg��σ��/��:6 �e�U���s �_}CK�:�MZ���ÈB�T�lq5s�m�y4����� �42��h3;/��]�!��%Q�%U>a]���R��UQ�M�[l�9f�`�dJ1�X�;|�=��#�q�^����6�p�D:,P���� ���?������Pt��g81���3z����0^2��`9��EB��fSn�Ґ�:
 ���U�`�����M�'���"�赨!��\����{k�O�U�����x���ト�5�*�-�r64M�5�����$�8ۧ�7�����g��5 �X[n{OL�R.^,��qR��AN���H�Cu�m�l0�ZQu��۾(�B5��!"�U�z���<����XYA,���UI��Os_����b t }�*Z�$AX�Ǟ0s\��
���1���؜~�D鏠��"�Hm*/,l5�-b����!뵠D<a�����'�/=��b���6�9�;�ښI^�ߑ���_���{��q�.��[/�w����*�����s�܄+2Dj(��B��%#O�h����V4�N�����,�͟NJq�`�T�_�
���t�F��q'.�Zw�No$���5�"l�Z/}H�Ix��#�m�|xQ�#�G�H�~Ī����b�r8G%TK�Y�ET\�2�`��\\�4;^�unC�X�3�2{�)	�S�w���S�Јgu�`�e�V��T�f���с��q\�AF�k,�v�@Q_��:�ULrC�%���W��Eq��3�fv�O&G0�-��r�|�b��>�\��e��h��e�wl��9�E~�َf�_�+���� ���}KBG���_�kgP5�h �^�n~
'�� 4����e2����Ӝw�K]����$e�N%K�?D�l��n �a@-��Y3����<�?����2��ܞ�rF���8\:�5�J�%�o�jݹZ
K�ϡ����;�s�(
z����u��S�Rs�Vi���e��������%���(�$W��f�K��
/�/�t g���v��۲����_/"��r�g�gf�^�" �35�[>?i�:���l�е�T'���N���D�66��]���dvA49��@QX�����,���?E��L;�Ƃ(���s.蒙�����{�*c4W�!�bt�9�#��� d\����J�y����P2"dMv9iBg%(9id�5M��ʛ��xR�w�OAi�,��
OO&�w�>n��}j���4r/��0#��n���+O踷�p��|���RO0�������:!�f#��+��i5iK��c$�-��+�j�4⾡i��^?���M��g���q����^~�J�O�j�[��(V�ݜTGP����=�|eY󙮏#�B����(��:��X��: �I����9�?*��44�D�|'a������T�K/]Ģ�kd<ǗRs2����m_���b����ذ�J ���%ft��@p�����鯿w�V�ϫ�	͸|�}0"p�3�u�� e����M������}��O���ID��\���F�-�Iמ�ggF�u=�\W����W���9s1n�y̸G8���̊���_���ɻԹ����=+7�Vr����< �XY��~R)õ�M!p�X�A���QA��p�����ra���*%L�u'϶?����8��"�.�i�EGl�2�/I.�	�c=|�v�?�|U�G;5����B^��Jy�v�&,Y-Yq�P�l�rQ=��p�Y:��\>�z�.:�j��q远J�]��-3+��2J�����ӯ��3���z���B�;V��V�l	1�me'S� ��ۧ�t�����Y}��/5��5*j�xGtiV�_cp�ko���:=
��/����Vd?��n/D�p����f��&#n\����M�⃉�* R�qA����l�L�^�%cL�P$���%@,��Փk�#d"�Us��3c��r.!��M��\"�U.���C*�����d��s���A-.@��k�ƒ��?�_6w>�2����ZX� 5��e-����5|�wX������[��O(<���O�*�m�ȼ�����'����|�)�u|���@���f���B��aV���I����\���\�P���_KY̪� 4��O����]=e�?�Lu�_GT�ok���4��:�M|n��R�h�w7+l�`��u�{ǅ������O3,��'ֽ>ѓly?*����{A(Z� �j���j�~������I�D"��[+6�� �GO�U�lc���#ŝ��ڐތ.ٜ�:k
���OP���hb!¡n�@�yZ��c�i<�H�p�H?p���\�s̞����s�"�y�t�#<��m"�]��䭖�'.qпz^�+��B[s�|reV�8ʹ;zX�]+X(��՞�q�T[.�Fz'N��$�r��Y��l`v��޾���^>���S�b�N�,gQ7zWe��O޼@FE>	�\l%���d)?9������M*��q�8P@��XJ:�N|q�J�`D����:��{���`{�IlM
-�䎃��d���F��o��kOt���s�Q�_�\F]
�)o.K׮�}�|U��\����*�Wh�v-S��NY��(UeO�aWk)Ң0F�_��\�h����Ħ1��
},v�3XG����3=-��W���	E��F�8s����cI@����Fa���2U��ۂ>B�oyٸM	?���-�2�y�;'0��u�#��rM�D���B�ǔLY�P�vd�����@�t�j��S�rB�s�o�!]�vj�R΃E ��|�p�r���LQ�.���kk���������[����進5b�.���"���g�5������ hl���c?�G���4dH��{ɐ��4]�$������ ���v�q�%��f{!��b��2�C�`���AHlQ��Np�g��O���>���.�Ï�Ck�΢�x�u���I�Y�N��ܦ�L�����5����(tށ+�ks]���r�6����b�Z�I�*.�G��e/��A ��+Mz��(ʫ��.���2a�$��_�~	���[�D���ǩ�%����1D���A7���*�>��֙X��ҏzu��D�L�e���<=@��R��g�~�na�<��<;p���y�ɍ��a��-]_����a�ۚ-�m��{������	�)g����,x����l��_oՊ��1a쭡1�b�����^�V��!��j��P9@�| ���.��_ XiU�3�9���0BBCm��=�8������g|!��w����xf��Sb�A]��P�_j�-���K���f{BX�d�}�8��9!�DJ�&�)����VF�2S�GK��;���a��rK��UE�~��X��xCa,�54�L�T(�3�
-ә���o�՞����Mʙ�T6E��2��-��5���6M�&1������((�g�}Ȥ�q��0���%����Cg��o�T3�Pb7��p8���Mue,��C��	icC<�s5~6(���$	Q��_h���Q�6�ߚ�4-]I@�W�Xi(�'�̠�dK��N���jb��|��/�_	�s��9yB��pE֧��%�5z����Zd�a(-��(�:]�wg�EaJA�b�Ko�
D��^,V6;�5�|f_�\T�S�TA��]��$�xGG��d���%��y��K�n�mͨؚ3����Hæ�{������3
����Qa��)��qvI+wv�-)ա��_���)[ ��\flR(��(ؐa�o^cRI�/2]�;0��|	q��hT�6J�վn�q0P
��v�]?l~���L���AU~o?
�7�HBr��t�_s�e��Zd�𹮁D�������k�ϼپ��f�+=��X㱧�p��r�� � 0Uψs������#u<Pk�U,���z�&��1.�4���'�C�����S��	.
Z��_��M��\�}a��d�fI�?�EY>���um(�'� ����$��[T��0 �R����Dxv��tWIs�@N-�1~��1<I[罂I5��<C ���I=�Α�z�}�����F�-1�V�r�K ӵG�[�;�~�{��Wm0���;pInu�V6x	��jl�^�/��hu-[������
�j?r�(�)}��(ȡ��Y����� پ�qk���S�]��$/X����Oy�(q2#���e���c��R�wc'T�Tۏ���Y�T��0�3�\V<�^ ����h����^q��>�yO}&>������Y����&�>�m��� ]\F�-Y@��'NV����b��M��+
�lAv8�iɐ�o(f�#q�@�(�n\9~���T�s�T����c߁��Q(�=o�M�|���� �$$î��	��{��u^Gh�,'ō�����F�5F8���o�W��$}�Jd�y�n�b�����1�rѻww��z��W;o'�@IC�#m��y����,�z� �U�z�/r�bʷ�aSd�	:W�,H� =��e���Z�<
��׼9Ų�#y1ҝ�=wP)�IzYS�@�{�)�/�7��؃���R鱤g6��&��Χ,n�+R$Y>�7��E'�˖_�6 �Z��٥⎖�u��?w��u�t��ȴ<gMj��;�!�iK��oߠ>O��/g���k���5iĞ=cO�& ��8�x
��A)�����y����"ɤ�E�
JU����w~Ҁp�2\@q7>��^5zyʰ�A������}�7�"��K��E��*(�4�� ���-���)Tc4��w���Ԁp�3�N�4�L�Ǻ~�q�{�bl������H���4T�9�u��m�v ��:�\ly�\ތ�����������*­zT�Lq�	7�/�C�+�@�?P��CA]U����MT��h���%��@m�.��oI�1jO�0s:h*B�a7��Ջg�</N̗TJ��?/S!V ��ȑ�\�ȃ�^ض�0���2Q:�y`[��0�vkl���Xʹ��N�K�o�(Jڷ�[��<=U��l+��C�&ո醎pB%�Џ�^؎��.,0V��.5&/���s���F[1�Ow�E SMh66�C����UJ�>pՉ���;����q���"�������a�Q�ٴ��B�.�rZ�v����ǐ�I_���}H.�Z���礐�aT��5���G��0d%j(��!��G�j3��	D�r�Ֆ��Nk��R9�e�+0�-؛5]�&�͏ +�qm�:�'�[6>s����{��^a���
����#*���{�B��+T>��Hos\u8)7�*�oC�d|3�h@����r.��ʤǖ���旇�� ���n�r�e����/���x�ի̤CJ��	��l&Xb��V����h��8�Ɖo==1��.����z�4}��jL%��H�n:!�����i��N��J��e����עP�ݍ;a�"�لnL���>�
b�|�ȯv��{����e�+j����Πg;���p0@�b�����of�Lk�f֌�E	�6A���<��֯�Ω	PQ��(:
��$�ߘ�ޠ�f�>a�
�?*V�T���q2^j�t���_,	b�[�Gz���dP�z����l�����Te�(��������K)
d��6�+�Ag�q�
��фi���-B���w��uȤ����ȓ���i�s4_y���*"�_�+�9����&L�L����4s�r�F�3q�ү�O�b]]U�����~�F�P�٘4�4P�q��Xv�W���-a�g�����
�W����U�˲�8�Yl�#ڨV%5�\��u74�ss�u�C�������<$@r�P�&f?��[��C��m�,�g��"^�K,q��O��l��O����p%��.jk>������"��T�������L�mn��堎�n8w���Dő�6���Dx�n{�Ō�KR�"!'[���*FL;2BD�l�֣�g�z�9�?�����sv[[an�� Z\����zd����v��b5Ƃ�Q�ӧl&Uص$�މ�R�;-�3�K���pp�z��"8�Z�us��˔�g�3�AQDT�Ol�x
���J5��Na���/?�@�x���Nh)�˝+���XE$�;�����5ޯ�]��x��vr|\�cԉ�Y
�zK��#H&��),��9���y�#������x��[������^⣣��h	��
�����	ޑ��g��NC��_lmд��ᝍ^�,6bܳ������J�+m$pih��A�٭�{F��+n���ì\N�z��zwX�h*h倣��c��^w&���֟vO��ź����7��CFX1ӂ���9����e'���������sRA�܎D���J�5Mtܷ��J% ��y���3���Ȗ����g��yl��p�S�o����7�mą�nBW����c�S�oI'�C��+י㙵3`��|�^����w����F'-{�_�wХ��:�s���L(�h?)L���dwUbq���ADj:|��7L��Jmc��Y�T�'�{�{~��Η�y�o�}�w�3�a<��F��炨֟S���u�軠���D�u:Փ��%SC|p�_�9��r1��>��9]ɍuM{���% ������4
W��ϹVZԌ���h�qY��Dǧ���-���GlZM9�a���W��H�ZL�l�.���llQ$H4�KHvi�ڶ0�|�Op=�N���+ڃ:)&h3w��/u�w��k�A��)��(	ъѦ�JK0-Ѷ�C��ߛo�)O�1���]����;ua�=mB�&��/�B��'ĿT���=(}�~!ٟն}r�P0k���B��Ve5ŬM)��^xr�w�s2����MXb�+�W�6aNX�$�<�zY�>�'HKn�U��	�2EJC��{3
�еdC�������N���f��:��(�-0�=Ω'u�E���.0�3�H|�%#��1c�u
���C7T{�	2O�a�s�lvzp� 	\�P4й�i� ����Q� ��ա�v ���˦�����)��ɾ�k8�)9� ��6��إ$7fn�ur���&�.�G�S��܃bH��9ԐV��/^��)�/�� t�~L�o�f��p$9{�MM�Yu�_S*�M��6}xҴ��@�
���Ĺ%J1$`v	��ƭ*0����L���V�dD��"�+��g���h��U�eA��X��OsF���λ����m�Mƶ��ڢ�UA�]���e�	)�5/�����?t1*���F5y�t��ڒm�Γ�����Ϥ�0X�2�-w�{F��ـE��B?"益��7�FLl"��G��T(B��b��*F�:��>�Ǡ�kz�Q�����<�/��W�����1v�0�O�ڑ���!�>Ѷ��A���k(�	����2����$;�f��$�ȗ׷h��F����Df��ݦ��V�q{l`�*K'��r���� hLsԈڞ��P}W��6-8y˴tH�fg뜅j��諓cdU��(�Qh#� ���p��6d#�KB~�x�f�#*�
��M\})���rjW�)����Ģ<��=�|�����Oz�� �����#+8W�E�͗MߢU&�N��������e�����Y���a)wb�����N���7@*��I�ukP� �tjD��#M�7<<9k���M�9�r�:3�j�N�:�+L��~��mɱ��L�IY>�����!��p�E`�� A�Now���������0=��I������06����S�3n�{X�0����� �7��5�v;��:�����؆J@Z��_#}�۸:�f�.�Mu��bc�3xPt�dU�]ć9��O���nK���oD��`�P�콀�����9�Y3�z�K�����qL*\BJ%%�U�o�oSL�Z��x1j��s�'�<w��%(uZri�����̌�]En.��9%Q�m�S�<�{T*����Iq�#g	�_<�"�ؤ�$���.�����\������ 6�p��R�α�F��3�:�U�5@EN�lPH�!�I��5Q�s·{/�Mh-�i�r/�}�G�i��[u���m��?a�;
��Oƛ��� ����Z=�ԡ��0M6��&a^���l��u��ϔ��<��N(��Nv��9#|�x!��*j�S0>hz6DnH���u�&��*+D��N����n��u;�Xx~�~Q_�i�c.�ɸ�M�p�}c����}�M@:p��������CUCn��'{��7!��*��Z���Co���R?������[������i�l��6+-?��󸡅8?B�=��W�q��g�������%^��"���ֱ�c�1(ᓻ����k�$i���ue@���R@����}�&�o����TZ�f;|��0�jiRk�>��@�$Rp�lQ0�0'5�	��S3�T���c�I`l�{j�#�F��3Z�<Zϥ9���4��{�b��Z���j䒒��Tv����^�����d*�9Mt��.l��3�M(�}���j���+P���d-�$G`�m�~Y_'����;�o��{�[o���%n�vo����[{�gL`U^�a�?;��ͯ���]�I��EIҧkȂO��t�>`8�IxOzJz�9��<Q�Y�E��~E 3�����B�j�a�Xy>�>�����mh���0�,�"���3�#d��l�cxW�h���U)c��ˑ�0��V���\�ʓ�aL��	����W0�42�r�P�]�.�ʕ�-��àEX|��`B������Y�]�V�w��]	��sC���.3��
-���_m�)�� �y��JS��عY!"�E�x��m��;®�e���ogiכ4�[�i�f��( ������V>�x��	w��0T4���K) }6k�X%�%�q�S����#_�-Ѿ�zt����G,��lΒ-B,�0 �㞐��6�8�8~3d�'�K�D��f~In��k){�8������v]n�.����L��Q����B�]q��	�,��r���;�U�^�C��Nr�H�_��|�"/��2JM=p�J���|��YZ�<מ.2�U�=iX��~��6
w�@�S�.�Hִ ��#ZM��z7�
/C�R�oB�߻�������^�,M}Ռ�T3A��J����V���Hx,S���4��f��av\��_IM,j��]�z�ٚdۍ�(&��y�a�[Fa�lڥ��v�4>��]��~�v��L��_�ᬨt�s��9Lq��lmA��ΖA?n�1a���Ct��*t$8�o?˴,�U�v�d�,�pf��o�����s
�*�x5`��S����JO�#��%^֟-ә?�I+�]�g���c��D3��N������j�
�?ȸ�Q�|/r��[�����!o�E����V/?:*@�SL�])�m��o$T��U���F\;["6��7����� |�Yl�P�g;}�8��O����J*-Fi���ව��RĶ��u�����`�Ze������T]�jX{*����aȧ�>ܘ��me��"�^,%��C��-}onu]{_����8_eQ�\~{��nk�a�ΰ�.��� ʻbEO���U�o�;���N!He�8B�V���]�L�����c�}1�Uc���萗�P��$ɔ���r��B�˷�ƨ��T���+��^�F��/����>Y�;D��\�ӽX��Y�}٠W׾�}U��+F����c��C���pޘ?�kB	������`��Ud7u����i�nh/k���`�		LD�WB#�C�5�c� �(�������ܬ�9���̾�;�lE�M ���7Bnt�y�esy(a�hԮ�R��^��#�gq��v٪���yΝ���N�9<��A��yc2p�#묎b�|;}:%������	�=�ξo���~��+%��А"��k"ش�x�N�	Q-��4��v�ȭP��#�J�Xm�w���W+!���*�HҼ��~2��}�qFr���kU��`�hU�=y����^  &m�@-�J.S�e�u���t�5�<�#���R��>t�R׀�z0���jU�Ԫ|����F��P�>��r�g�YCƝ#�dK�()�����HJ��0��6��9K�e�ɚ�$������F N��T�7�<��$Q�׆(@��w.�I�#�H�K��aB�M�b{�p(�]���a��NBW7T��V˰^����U��a�B5E�彬�5}?@-��T�̨���b� ��åxg\�I&6��Ǣh��Y�Yw�ݎSXVn�: FQ�9���i
��n�! �ї�o%��1)��K!O��Ȯ��]���x�`�ss{��JiG0�J�ݭ@��y�iQ$iǌ۶����Y��LZ\fE*�?h�L����,�	0����Lx�:*��Q�!vr��T$a�X�aS;u�dϬTl���E��#�lN��[�[��O�6�q�U��8���gH1n��P� �3��ua6���-��𴬟�H��5s�L0݄5��5R���=��\�w�qg��I������ ��ǟMԢ��s��. "�D�4x��g�I�]�i^�J�5�t��Y�$����,Լ��X�MY&���4%`��T���Hdt5�͕�ҤB��_��< �VUZz�� �x���TҶU�uN�mh��� ��!��X��O!����oSfq^��N�vD�C��o�&�)Ś�{������9����j�%t��n]|>��� ��8��bT�l[�:b��#o��t� 5k�����e�Xr��x���e�k-����z*�����/�`�#S�����<{p�K\pmL�-�瞡�R/N�cr�~�O�����kIU�n��`�o�2a�������,�q2�)@��o�|]dW슲\���`U�
�d�Qv����{��o^�:��kӉ�m5�"i��\/�u���^�]�y��/��Z�ԛ��5�3��Sc�Y�K�q6[�4�}�]�-K����"'(\����M��1�7��¤Z��`������k���,��Y���g�,�"�ħ��kSևd����=�������H���$��n ����\Z}���<lH�c�=!�.��g뽜M'?@�����s�G�zg�X8�n�=��B���J<�s72�6����y1��yCAݦr-��?�J!rX�������z$qZ������٫ѣ���t@�cT#�.K#i�a���B,�n��(i��9P���%<f��X���W8��q�G��PS���9~"-YGhO���'���g~��%>�icg[�����?6^Y2�����
�g{m��d�>-GǙn��y��y2�)X�}J�ٲ�<��h��/M�Ex���|�D�h�L���O��E�����.	����Y���-�$u��I�ބ2qD'7lD;��h��K�����@����zj<$�pT 7]�mɧU����qc��/�;�2�j���At��q�Y@$����Ӌ6)��M�T���+4t��
�j	�-��q,|���e;�j�'����U�d��+S_
0aF�
����T�<����UR�r��&pa.�}��a),�(?�J��M��vY���u�C�1��"|���]Cm��a�tHՅ��9H�c��r��~	8H��|�$Ҧ�-}�V"b.�o]"_��L�P� s��͓)�c?�7f�@1rZ_�*{��������K��A먗1���(���������� 0^X��9�3k@�c5~�&���+~����$��k�䝀��k�M�M	��$t]WC�]���z/l�#�dbԈ֑R���g�>|��%����O���%
u�r�kP����o�r�;Wg(\��H��+HVK���ޯ@&�� U�������g��rbmǽ�&����z�מ������^f�9fX�CO��3a�U%s�{�ɐ9m�����l�|n>
���zEc:h��k�����'���j�vNPBkiTU;L���t�*�{�3�1�����`��g�\�B��O�D�#���ߓ��S|��+k���3��4ub�,��1�+V�IxV��2ߩ_�K�~��i��Qa��I��c׊r�d���B�F���:����[�����X�u�2di�if'�����Ɯ1�bp"xcY�.��r{���4�����k��Tsb�>�֩*z��FN�̟8��E}��˶�9ހ��E[uЈR�%qA���������g�ٗ/ws�qM�.�A��(���~`
�b0��0��b����),�H���\�?>R�k��"�a���I�ʴP~+�8�)	pm�H^D5����A��$��=��5��׀��P�yj�4�y@�Ԥ�n>��(Tڊ�����:�2GL�ڞ]�i�q�^"G��y���$�ZH�*��o��/�yE�@������V�NA|�K��l!�L�����Z���C�/�t�������|�YN!�c�Ekl�˳�:у=����2|�=����j��׮M�z=g�
ة�Dp��I�~y���2��ۻ�8G�N��[�D݇���{�D�,�2�� :�6�T-��*�P5�/�Jy����ck�)����0���y��\�
���M��]�,�vM�pDX�].Ka����w-���Ml��!�ȁ҈�=&~4�$C��<0��_3�+]���-�>0��GFw���ϭ�[�*�F�T� ������Ll4��<�8��B��zu6&�������O.Td���� �?�nߍ	w]{�� P�l'y@ޕ�f{$cR������K��t'j~����4,�R����+E7p�o������ҷwiXq�27��s�a�ZILp����m[�R��#F��R��;���r$��-��e�j
���@�C'�`���uLgGmJJ�JY�Ɇ���T�v)7���*���95+��:���m��ذ
J�������0W#��T��;�c��c���k��1�&nH6��BVB��F�b˄�<�о�B���L\]������J;�E7�St^\��.���]ָ��n'�+����ݩi�=qR`���d���������%l)�8Ӄ
=��#!hd���Yu�:�1Y4�ø'�<�2{糧��Yn4D�P��\���P�6����d ����οi�q��!�b�cy�U�)4�%��M	�_�3G��l��,���ddʕ�=�XZ�SG���U��7+|�'���Q��*��?�2�C���9Q��(�X�	
wl*���ӊC���I>�(a�P��-4q�[^�I��%����|�ڛ�6D��\�D�IK������rY��̵��C�S�5a�_�����=�&��y���C�q������j����f����
(�J���D[�S�y���UbQ��z&��M����kG�}���z�RAu5^*�Ș�l���l�"`a8F��Q�V���n�� (_ �="��N����dOXC8��J�a	,a����n�8kuǁ<��"4��'��/J�:0tL5��H2��T������;�2fh`�d(��dI���k+J�$8Ɨë��P9���nifYC[>~S7��Bp�"���	�0 ��*��Rd	�l�@�;X��/��&='�w��z�P��v���?e�+��S�m�: (�9Xs�����u��nݣ��Nѹ
��:6�5Ӄ�B��m��~S�(�ELs#��O F����m3�v��e��u4�#O�kMW � �[��v-y��wuhJ���6
H#�T3��z�=.�2���%����ƭXgU�g�ݏ ��B�^�@�z@��׍�d�<���q���v�dV=�l�r�y[�Y�xk |v�k�#�k2��A9��*�/G[^V�{�	�S!�� ��{��m!dm����� �|v �jщq�"",�q������}�ۍN{���~M��!���}�%�4�U*��	K�]�9��M��ݫ	���Ӗ����*�Lo���g�}!n��@rx�*�n��i�W�G�%��p��XR���i����3�9�`Ƽ`;�f��4w�g���CCI��+4{��4��X,� Ś�ہ�)_�)a�@kcC���<�97#���4M��\���z����RyeO�̆p(J}1��;G�M��[�(�"���{�O�	!��<mj�?�*�<����=]/lFZ�T�-I#h��p7��� �6����m�b��)�<���Q�/5�@Ӊ�M�+�($:�;����]QI��R�((��t�?N;
	���P���?�����J���]���z�YaU$h���P�=�d��p�z <��1�x��Źq�xap��4b��1nR��2��;�,~��Z��N�4tՌ-0O���:�ڑԧus$�t�4�5;#�Q�\%��i7A�Jr���Sq��*�yzr]�R&�����aHں�����$)J�ۢ^������3�� ��Y6�Ŵ���ݴJ㓲Q���3������=�Q��JC�v�Ԡ\w}J��_��ʃ�����ĸ.�Pm/�Yp�hrd��ڬⶲ#�Ò{��,
vU�l����e/�Z�����Y�e(�O��S��q�%��me�2�#6�����.�t�Wo���1��.�q�
�ű�}d�(�������1���*��i/'�$�×tK�0h�$#!~Mf�,��ad�w|h�7��''��O���.�Ynۛ�|�	��ToM�>����!���a�6��9}�h#��T����<R�(U�FT�3��K�x�e��Iy��QI�c�D*�E)�uo��]����.���c�A�7��}w`�-�r�Ԃ��ٽ9Ag*��uU�rRiۄ����tb�lT%��\�n�����r�� NI1�y���JU{�� w�M�Cd^/8B�s�Mf�N��Q�*u{I:��f͡��(�a��|O.��{�D(��Fp�<��F��+^7��r�ju~�aq�M�(�����8�w|X[C�O�5���6���-F�>M�Y��w!�������������)/��E=th��I�Is姶޻o7>B��uqc�|� y\Q�(uٖ���D2/p�����w';�*�.w^1�<����[e� �0�o�:gF�1қ�D��3ף�����5�6|��4G��'WbK��Ɓ�z���([�+?5~7�j�!�~��M�eûQ\3U��{��K��v���LxL���B�u�`��t�ի����.���MZX���?�e�4�� ��P[��պ�l?j]�3',LQQr��	ly���0���h1\���n;1t�u}*�"���*�B�4D����E�_qŬ��k���Z*޸q�:e���ܑ��Rz|v��K�ɸH	.韏�q��b�+����.Ra��� ΁fq��y5�J��Ҿs��x�r{�ч��WYyy6���k�'��V���K�N^�+J��|1�65<���s�AMGO��![�[5B�/����"QΥ��Ʃ\�����9��tj5��B�t�r��ٿ#D6�v�0�d�ZAoمY�thb��)}��C��7͚�����!&�&�5|��9|���lP��C�o���{j9H�����7����j�r׸��C�3�J��(PK7u��O���5�6*�T� �ϴ"B�j@̝fɀv���Y���9��uQ�Viw��C��=e�޿�G��=J�8�	�)l�F�5��l1�~I�o4ѐd6(ōu��E�1B��?��}D�-�u:��d�ve�����l���<i�^����hL֖�D7�5�{O"�n���>����__W��n\��$�0��62�B��:�?�yj�.O��jǇPEy�b��Z��[�0�Jm+N�F�^ٕF�W~+K�f�Sb~*
��J`~���s����vg`��MG��V��C���0
 �����-N���:ľ|��J�Ab����I[��� %���~�X��>���:XlB�qXO�n�<�2!F������h����x a����G��VF��e����t�W����H��8��L�Цz��/��v
���r���=#U;C�3���!Lչ�郾����$��\*h6�.�c��������fn��`.P�$�9w6'���k�3ꡉ�t[����C~�N'^��y��������0Z�0:���d^}�\Q�Q7�CfASo���?�u�b򶗯�{�Ro��4�[c�݈Ͱ����5"�sϔD�O���kz�D/68_�����j_r�s[J@����q�5�x!��ADsȮ�x���Ug���7o� z���ⳁѣ0��Z���)�B�&X[x�w[��q�U�`�*1�ś��8w�`$��/�)k��|#4��E�}Z�o���Q�/�1)>E�9 �\cg���|?D&��)_hzKZ0
a���[+-�9ڏ����I[C*��I~��,��I�Hr�� �D�8��z�r'�L̠v_���5��I�&�3vj'�Tߧ����4%a~�����a�����D��*��i*�/0���)s@%�"r S��+���d�z>��N=�{��O�󦡴��-4��v�.�mѽ 5o��Af�����f �,�������$���#�Z! ("�Ю	Y�m��eZ��</��d���B�gO�l7�o�p�H�tE0+���D*�]I����C�d�q�-����{H)��#
q/3{?���MÓN�����N� �=!�.-�$Ǧ^w+l	7�����U�n�E!k�����+>'ǰ��K��}?�Q�SI�/"׵��H��0KS�Ѭ}¬��uV�1�oaF�-�!�x]˵�*0]���~.��XLJ��+���1�\�S��J���-aaZ]fI�xˆx�� �q��O��F�I�E��3/%,�N|m�<�U��-��7���Rµ�i�-q�?; F��t���e�9?e�K�C�}s���qv�:�wPeް��b�r�q�����=�c�?0w0<�ߥRa�m~��.�_�-/�$aokr�Lyc����h�7��n��k���'5z���n��u��9W��	�d����g<��sȺ��4�#�����f��즲l�	 ��]�֨��	�g�۩+ܺ�[����C"��(��_��0V�V�Y�$�Z /v��k�4Tx��|l8Ҹx}��O!��=ZH{㑨<��X��([���=M�+�����<V�TsH��Ҙom�A�l�7˴��ρ �hZu�]7cO&���W�4�U�
�Eb�si�t���\����+v�g�Yk���
T�~��ޢ�xMp����Z��SьP�:]��e�V�aE�zefh�qV?�7�^A��E��.%���;Ǌp��b� �茪0���nM�Do�C�JLi�JD��z:�Ź����v�s��_��'j� �L��'i��t��G ���O;�G��IC��&,�j<��|g(5�l�o���s7��m
ݽ����K��a~���� 'KGI��E��Vt�0�UU�GL��{t�Ι�3c�l����sM`Yk�Zl�˧V���$��|���.���p����3g� ���J�\<f:V����c�}�ZSI���rd�mk��M<�{/ҏ��CN��j��ڠw�K�����63��Z	�ϐ��:��:RAV�H����l?e+�O����H$R�W�ΰ�dB.^ʇ�W��ӭ�a0mj������D��k�B:!�y/�0|�vV�({��R��TRSc��B��r�Gk�uF�k��w����(#�= �*i'�9֏��D��1|T*����� <��E����vTwbA���d��|�E��)+q�$c5IKH]����v~��?Ԥ���!/�|�k�4э��^q�ǯ�;�����Ydh�z�˹��/��+gI+�<�BS����_SgPY��6��>h@x 15����t�*!����1�g���._xt4��2�)^ObR��$�:��}5��)�e�1;��h�!էޏ���N+�?�x<x�UC2][X	�`W�E.��!�$,�1t���m*�YHC
�
W�h6>^����*�}&���`��6�4
q����g�tό���Ud.n$)�w5�Y��q������C__f7��z�8w��1���-���%q}	�xi��jZ��3�����ek�䰦�t�[ZɊ<qm��A\����3`�� �H%ǅ�|H�t$�؇�|]�������L����w���Tz�%`�,8��,>,�=�� ���N鸰yZ'�d%Pe;g��n����*�'�P�A�ؑ[�H�&�������*pK77�Z?J�އ�F��&�{��D���}�.K�B��	y.;�z8���g�sK��8��
���A�(xjy�����j��І����A�25`�0�k��5�W��Bڞ�<ѵ��Cv���.���0'��XL��\&����s~?� �>��@�
�%ۿY(V!"��+�.�qHjo}��,r���Ã�Y�-K��$%��"����o��1���<~�������m���@�1T\� �0��IR��p{5��I0I�n�"2�v��:$Kg�D��K�+8��?�VwY�b
)�$���QO)LM�7�"�¼cQ�5���Ï�l5�����ĕ}T��m�99��A����o�ps���T#�
K26��|Qx��w���q2����:t���u��V}j/���r^�m�ulQ���O�����|8��ZZь������S0:]������~�!���) f��D�N����D4����Bxҁ?Ƥ]���F���Eb�\����K�Ǒ�A���PFD���V|Gl�	��֨�3V~��h���[�9i����#y�ı�{���$An����N���jo�����T�W����5N���䠗�8���A��HMj�`]�:d�$�1I{���L�!�xe�)��>RL;�W:͋�ڒk%/	�&��7�CoĲ��c��j�g���-�I4��0��4G (q����gj��FV��j��-�����0�	4ܳ�4���#��@����Q<;��B�'��A������UlfHU=���3	VH�@Hus���S�&}�1@З�3��+,��HW��WF0�|2���̨V�p�t=t���cݝ$�le��9�4<���=����Q4�����p�x��wx3��x�m���9۱�~Ec�U�T��Ù�"��K�(�<������[�HZ��>3�:蛃�)�uv��p^��ƷODY�6Vߠ�{�D�������O���t�3�:���';��V�oOR$�`o抶Ph'����*���aW��s�Q�;\fK�3(Kٴ���i;�8��������a�M��iC�b���$��h�����
c������|�����x���60�R�r��B3�mH@lk���t�Gz8���]�{
&�eD�r+��H_0���}t��4�4N�#-sk�@x��=���]�a-�Un/m�"�~6a�Q�P��|��]Y�;��'ɽ���ee���B������`w�(��Ҫ)���ъ*k6lc<�h�ћk���������xhmX���W_�]� ���s|'j{n�Y����B`�����*
Fiޛ/��T&&�1����M�.LF<�1��A���0a�^S�Z�1*��x���	f%;1�QBI4�-X}7u��*'��������8&����"������~�pA��qg{~����!^й����潓���h1a�1�o�k^�C���E��1����_̑\m7�(�&bv��E*�Pt|���5�<�|j�O�P+nLA�az�@d����n����3��j�F�{Δ��b�ed�63����}�>$Z�����|�� ��"<rCgaZc�v����WH��~Y�y��])� )L=в�F�������߿9w��!+X�oT����4m�
E;�Ն��������d�Y�F?�C��6J��eua;��3��<�7����M�m(^S#��!��s�t0���ɛ�|�<qZ�_�8�\��v\$_q���R��,��:��m��8\��`���9kU��])uO8+��y&�]T����B<jR�QcRW.D���֜Q��3���o ��^N�(�)�{�ʄ	�0����u���:%��C�:�l��̧]�(�����L3D��F��zP��W�{��ѫ��$ժ��N'��I���ys�i���r�<�������dG�{:
�<V��,�;"0�ML��_����� 鲥W��K�G�i���>RI#��w��!�*n�����/M���1��7�p%�Ƞ� u��zqeJ(M@�s��k�䖠1�W4A#�H��!?5X�^����ג�&���&hV]{����nv8�G�Ǆ�<�j�.��R+h1���f�h\����Y�������3���>��\���D���`�����������fF��L��/jDK1�0��������H�S���>��PaQI��e�Ԏx&���MC�eF�ATßy����%�X�~c�44`�1>(@��ڴ�2�E��d�?V��z������I��ց�Y��=�|����U��yQ��-��<ȭ���O҇�=�4�����d�7�ңJ<r �AxނsǗwn��_=$�y���q����8p�W������x��(�H��Y��hC�J�[(~����*���I�E�D\1�u���'B�J6����bO��6-���I�D��F�R,�pG�� �*�Z�S��}^\�R*E�S�iK�'4^H��1�x�� ��q��%>��!��avPq�GeC�H�2NS��S-�ʴQ�/d���y���
KgU?��)YS���qE���agby���IP����И�t&��˄�w�w��U�š��dȌ�6�-����^ǎ#K�R$T,�&Ox����s�}�懕��E���5���	�r�q�5,�i���3KR��)�;���PƄ�Y��=���%��Ra�M�5ފlR�4<{��j���̬O>,�gM
�M�Z72��-aJu�E�Am튒GZu#�;73��a>��z�#���6�K�����h��f�~�/;w4X�������*y��v�c���n���Kg۫�� �I1?��x�����ؖ5T*%2�?C�r]�e���y<��'��)�H���s�j9r'MW��?�N� {��h!� �9�z �XU���pj����v�cJ�õ�m}�YC��bT����8
&�?2Z若�`�vp���(n��&���0C#q��s�El]Ak�硻6��l�t�%���" �������]Q3�s���df��8@�r�
��V���>�`)�җ�*��jy�&FB���L��q#�B)� iq����ːP�T?}d|o�ŋ�X,D��FD�wӇ���3�f.�ۘ���^0���V6dAw��ý��Ƨ'�(&����oS�\So��%nRQ�=�A3���Kƥρ�/�Kr���S�ʄTq�g(W�Ի7	؜��(��´~��&Ta�����!P�qz2��}7m�j^;$������`@|*��tt���<���p�`���k��۸��I������#���_^Ufh�Uz��I�x�d����I�<*8��3�~��6�\���+Z$@�
�Eʗi�rX���I9����^�lWt���P��Md�P�&_岂O�J��i�-Ƕ`æ�S�O���y���).�Δ�F�/�m�:��EY5���OF"˝AZ[�K���D��H���v?2Ό^�)$��,LU�똡	3��S/�fw�J��h��O �����c���\c0��ƃmqGj3E2�N�������zL�X���?qJu�f*��+�"���tFX�D����;J@���F�]?��p_E�0aIT��V�D���(+��zL��`�hy#s�|�EkU���b��`�]��Y�\�F	�6+VФ{��� ���<4΅���%�"Y�#N5B����7��y�V'��&SK��."T�V͈Y@b�=p6�Ӯ���Uxh���ݷ�����k�?s���̤�@�ӣ�-�e�]XqB���}T`J�y�2?l>ܥ�x��☞9�R�<����%�� %�|�AoVb�I˱�R�U-����76�8Q�ϣT�M���` `�*��� ��a�����r`��}��*sCT�����fj�p��b�?TTKэW�!��۝���Ha�w��D�!n����ҁ��Y1LU&�'ܚP�,;fB�G���P������hw]�,Y$b���9���JbT����?������z ]9ع�'�"b�6d��Õ��k�2�&5
��QB�יk��ː/�3����z�[�0�3Dy�̉+`�!������k��G62�6��������}:z�#��&b��ΰC/��\��Ǿc���pl�c�,T�YP)i�s��+��s��XN
 ���(X9�3��>%�{{��Ip�/ik[���bTn���[�^��ԩ]��w0�	"��K�~�2|�	�y�/(��g]��;�ùM�Cj\gv}2)ҮO&	�t��T�*� X�������p�Ŋ���1�Pr�!]$lI}�`�����i�,�����%���Gz����Y��db�4D�'�ONʉS�-��&�V�w���ֲ�O��\��5��hpQ��!H���,	�.�Z����g���Ǡ���	��o.���`�[��jҫ��C(x�'�t���*�(R��3
K�ί�[�b��'F���ʜf�{�1C��3<���%j�7$n���?n�U��u0�E���`�h�kHcP�����3�,�e��#���=E�����J�*0���V�|�8���F�c��d��\�X^5`1�Б�]5����:�����^�yi���B"�X`���
ۆг�s	����c���˩fU:x��'��mn7��z��c��a�	sY��{ǣ���R�y���:g�ꍜa�	F-c7��#���5�r���g������Կ��b3�\�-	d�M��4f7�1�������F9��~�\ 򤭚�^����k�	#�7��zVE�PÀI�Nn8�<ݧ׌���Z D���0�8c[�A��1�YB��A�~o�+��B�Yŀ�W�����p����
@ܵS�%��b.�nv���i��>� �����2|� ���+'�kF%{��$��2>�8og�t*�^���F����?4���*a���r�]�t�Y$�����a�������{<.K=x]�r,��3�]R�K%�.���1���;<��XJ�Z ]�.��~��%gB�.
�4���~��T�D���3i�Q����Fq(jF��O�~nQ���̺��K ��)�� ���Lf�(u@��"ɧŪ ��xV������~�L�޼�=�7���0f�\$β�.V�����2�1��{���
@���)AB^��{��^[ċ]vO��@�MC|Ǽ���x�c���o��o������e#*�e�.��o�q~uf �&8���"�Ɍ�́^��;��4̺�G�G���>v��ќ��o[x��@@�0@js�rJ��9���͓cܻ;V�O�b`�u.j��C���ND�*8�����>h�4_��x�x�$�ԣRa�?������)7kЍ�L�ɉ;.�T+�2�e�/��rȟ\#�f��#�fؙ.�r����&��3��bh�ǅ������\w99����}�4MOE����9R�c���Q*(�7�>#>h���.2"Oj���w%�~9�_��� ��Q!5pza[m�E���v |�qA]˱׬بn�~^U�]�����/�r�h_�;�: ���@���`����\��=�"�k��Q���&
:�{��H�x:w��ɻ���?ĭ�N��WW�wy��8��nQ�ՌW���b#�{^ɩ��E-rj���DX���~��+�u��`+��3�GdF
fC���\xG�`}v��Zg<;����׻���t[��nl�'�G"2%��;Aǿ�+ž�m��@�e&�=�ֹ����^I�փ�EG$o\=�`�l��o-�'ٳg�ی3^=�k8��K.vJv�e=U�gPjg�N�z�̃���U����h��шx	<�E�b�I0�2�^�̗�������;2�� �!#�qΨ3�Q�����V��~Nn�*Sy���Ԇ,�TJ!fO�.��h����/u��X���M����a�};0ިJbX��f7w���q����>�����H�+su��ɳ_xvU�s%7D��נy2�i��T2����'�x�+��ӽ�	���=��R��1�!�(����:�!5B_���-D�Lkr%�T��w;�,P�
?R�^6�Ҟ��.�g�`��؋W{g�rߑŴ_�D0���_3���|��;�-�A��j����(-���X��~��i.t[���
��-"Z�Ι�O�k㽲F[�3<��_�0��\YU�����d�N�|��6m�}�j
�J��:J���o<C�t3ܭw�;0��{w��&�y��vWb�5�_�'�����a�do.�[J������"�-��^i2�]�v�`.ߋ�S_hx�Q�m}��Ë[[m|)��HSݡ�.v�<����o�g��4����}9E�A*���pd�M�pI�;|u���Y�2�48E;�܉��{���@�Y�����k��$�#H�y$��XU�
� �@u�澀F.�B�����م�k�".�O��)��&Ry���+d`�9t�'��SG�-v�7�H��	�~$Xuu~�N�K�;����M|#7~hVq�o��׷�Ԯ��|�WE�h�sW�����SWո��N(���(���� qS�����E7Ok�/��͂���Ǳ��[q�O��|[�L��Ѐ�c|���~
�*_�� 5
Ù��{�%k���V�\o�����K�Ԗ9���rx+	��P���Kӂʞ�1G�sh����ى���V����Uo��z)��Ww_X�����A;!]!dJ �e��Y?d�5���vX0�l�qeD\���A����a�x�K���� �j ��f��.U�Vo���^,����B��h9��9��,?�`��"��sW�뀴��J��D܋�����*�9�Mu�f��ɕ�V���/�"�`��������#��ށr#h&�7A`�|�>�"�g�q��ei���Vh�S����F���	y�Wdb��F���"UJ���r�����K�f2Ϡ�5�%@	>�6P�ȼb�u�Ҍ)��S�z����m)&~�^�"�HS��L1�p�|(o�K�L�Y��������N6ŕqt��6����?�9v��W.�$��RZ��<�����'�'�-!?�Ƚ�ׄ4.L뭪�jBX���D�h��1��-��N��Q�f����#&�"@�$ݰ�Ȥ�W��]Kaf��'��"�����{Sp�Ճ����3���'�E����J�!��ix��im��k�f�g�f���a
�rz�ҕ_N�ЇC��L�6�k��4^�7[:���k�I m��zG&w]G^���ŦM��D߭p[�gma�����a����̊6�E��b����!�s���y,5�z�Y~�n+����Fi�lL��X>Y�R3�~�vk)�6��R�W�a�~㋦��� ��t��O��,g~��m�~М2~��ZyI��)e��E���(P"����#���p��|�E���d*�z��l����'.���Z��ǃ9�QpO�Ӗ���qo��G\��Wy����1��i ue�ݰ�{����W���0
(��>��*�'^[��S�3R���y/~O��!�Cwݓ@���H�$Q��TT���?�m�s�Ov�ԣ^�0�4��+c���肼�T��B�V���Y~)����b�.M�S`جǨ,�MxoA���@��k� 8���͕=�S������H[���Q]�`�8���5�b�t��� 6����8��ւ3����&O�?q��Γ�ّ��Q��Cj��1�8b�b��(�_a/���d��%�Ie��6�x���,��yA�#d* L����n��&U:����/���ʣN��pC�o�� �b�0�D3f�)��:�e�3��rvX�}�=�'ŷOyU��gwBS�A�U>hUo��oj��J��P�B6�)�����O�ִ��!iG����XK[�y� ���9R�Q�q/�{�\��q\1k຋�^� /٨n��(���'��]��T@ųf '�
���j|s~@�R���!���ε�v&�n9c�؃y�$�<?B��h/�G�Ybv�&
�����x���l�v�B���9��o;EH�V��Q�N�P��x"����_�7������<�lb��������[�?%@e*��/����|�.9i�\f`��Uc8�p!Ao`XR���1�0mfS����(�l0	��^Z�]NS���4b����v]X�JF���>J�(��?I��r{v�[-vO�d�a���<�$�2�E�\��h��k	/�U����G���� ��yx��$��A)R�LS�j�fc!�p�_($Z:���ҕͣ`�C�c���U"�U�cD0�"��^P{1~�<q��ڃ5��;(����,K��]�TuY(�lcj�cd(3��Q�To�kD����p3�&�Y��҂��2&�Ū�&����!��jcB��rGr"?��ܳ�R�R�:�&�Fӱ�lyY�?#B��{�OdY�+�2���*�i�Fc�N�f�����4��up��W�9��&�"�B:�?+x��So���i�͌bv��>OMH蠞��;C���AU����|=�ҒEq�S<H��Eu,��P(?HbR�������RU�}ny:���kC?�����
�;�=^W9���2:I�tF"H�s�9�x�lg����Xڮ��o�rǙlկ�`����PkE�l��skF{�;;���*&Z�6�Pe���	
�,af��;�"����`��1�_�24�vBN��m��(`y����|"��v��"}�9'r�N7KE6j�m�^1��~{̋~�f4g�*BT�Q���V���Wf>�Y���X�mI���g!�)���5b�ׯa;�)Oe	�v�i:�t2�u ���>�z�	G�-���N�����L ��TZD�6�}�T���z�JH���\J�ݭA���T���Z�R��פ�����W�З����ğ�ʷ�;K5E��B-��%�K9o���,W�oE6T5M���c�Y��+$�<Hٷ�qp���'T7�w$.<�W8�V�EnK�>J�-a%��^"�櫻Xb�� �T.�$j�����f��R�SX�f�T�T"��kx ߣ�`eZj��裐��4��}FҎ�F��| 	ֽW�I�
�Y��kH�H��ܜM�UB�o2�@�n�"�ʝ�cÛ�����O�?�A�~X@���ad_�Ҳ�Է�l�b�8¤H-Q���2~��0�,f�h�@�Nbq�_Q�F�L}LoL�S
�p��}�5��U�n<˿e�=������T$��%d�W�{OA���ߞx���dq��G���ȯ%��1���x׎��F��'O��k�k����cy�	�-�Z�ơ����t.����e�@���7[��2w�o��Í��E��x+[^���qV�G8H�.-EZ-j!�c
�����A��"`��ٍ�*fC㎖s��:SQ(��,~p����n�zUV�����#J2P���%b���1w�g��Cc��LH(�#���5��#	I]� ����l�4o����ˋ+�QR&���9�� 4wF�2����q6�����S�$����N>�Q,f�	�j�n�����l��"�e�2jv])��%��Z�
�.93�7�^���d�}H]q�2(��pD?�;h=��^4�)4��@FN�i'~'w�3���]Z�����G.�����cuo?(��]�f���e������w0=��'��Z%�H4���ؙ]���zT�Z� k�&c�N��	d�w����ɝ�n��DK�������x�<����i��<�G���C]��"KS��b[��8d��_?Lm�w~�!���v��HȽ9�f�M����Wj��B�����]o�-�4R]�B�e4M����&���&;5����RF�h�Zf�r��������ʟ�-�t�X4¼āT��J�	ryM��(����N��)9(E�p�#��|߼��O�j�__,��� :2�����Ǒ�ً�"�|�=1׵nw�fT��'�1�����o�W�S����9I1�a�R���L �b���ӟ��Ax!c��i�R�~�]<T$��DN�Z�:Wa9o�R�9RG(�S�G��L�z�"tK��?�^����8�^I~��C7Ҍ��p�b�����=zIj~��$�+�cTi�O���C"����S���Z�Rn�+3�I�Y��mT���t��"0��$2��Uƭ������|&G�Rq��wQf��r�p��ܝڂ��㕞�GtɎ�q��������mRC0��QJ�'��q5CA]�p�c�*���F㴼��}�@Mw�;�!W�RX�=�hY��r{�*�BL��=n��񷧗�عƚ���:�Ů�t=�uX>,��=i9��^L��vu(�⏜k?tW���1���2�$'�D᲋��R蜧:���ۢ*3s�H���v�c��E6�v�老º�8�WwИ8H��gj��\�8�����?�\�u!���W�9�)<��n��ǆ��=�l))�D(����+-O$�3�z���4*Ζj�24]�s^����&�4S׹��_�z+�؂U�ڈ��76]p_����̷�zM�h��b�*a��:���#P�U c��t(�v|i���-�o��~��0<��1����%Ot�I#+�>}�����HY�Y��K>L�eM��A�-c�?mf0"�_�#'V�b��B\���u��#Bkž�y��$@Ӊ�>��àB��G�}��E��:����4Q�-���o�Uӂ3Ձ�������nۢQN7�?�ϋPd�3��Hcg�r�>{�5#kUJ砪Cex^"R��N-\~�LZ�Ss����"A�[R/�C��Rߴ�����x�"��S9�����;���7��g*��x���P��4�l�R��eMg
����/W'05��X�Y�ʉ�R�/�������g�� h��� ^^ʾ)�����Xs{��3�	�}i�O��eF��[����6�萋�����(��(��n�3��#��rU�}Njm@[An5��@������y	��)�lV%�� ��n[����|��q�e�bֆ �5s׆i�.�5���na��`����o�Q��G�'U�;�v��e��T��P�#��`h�ʪRm�z�v�}5�W��p��9bQ�jᣆP�e=Q�׌���w,����lD��S�#����"0�o%aĖ�|�=��pk�Y�1?��]7��ŋ�Q�T,�,��%�ꪵSvL"c'�d�';�߯Y�&���T�>pEk�,��9_p����+��g�
6����Z,@��iC�u��y7��K�������gD^Ba��8�?Ư�����.��ּS>��O�>������2^�e0�4��_�v��׽�g=�7�g��I�'^�t��L�\Ҳz�.>
����٩�ٹ����>���I[�LÖg��uDh`!a�Ͻt\!H�-���p:D(�R.{�L�f|���6"%��n��vT�A�ԃ� �ى��#<�"�)��]���h�:�]q�^}[E�F����Ylȋ1G@62�#̂�$̦Iކ�m�|K��/+�'� �FރJC����W�A�o���/�q"Y%DQq��Z�ԣBڇ����� ��}I9��+!2_s�G?ae�<�O3�vn���U��:2{mf�J�,�<��|Pu���=��z(�P󠑘��}cO0����'��$�7r2,{Љ!�
���!i�5*.�6��;-V��)�t�*:�d��z�(����W�p)��;3�rAu|�}hy%h�@�-k�ǵ�κ�R�ܛ��kh�k����
�� ֧���T{ח���#EaD�->nE����}pO���ʹ�х+d ��Z��r��	vfb��!x ��O NB/W����V�];�����-+�$>�S�A(�n�1����?:1q0�x3��ծ1���k�m.w��ߟH!x�f�t��s���!�E5%����������mΦU4��9���Vt����C�y������(���f"�q}�Ҋ-Q4��&Kƃ�e(F���0�Qϫ����/A��9r,�Ts���U3�v�[H�慱hx�?���R���68���T�?�5�0�u*=J���ѣ͏[�X���>-���u��r˸o��Q�c�3��x�Jג0T����w�GOʪF��	mP��W{$�6W4�㥚1��� �^ӏ�e�X�˦oC؃��~x�;��y(������1#�	T������ݡ�s[�}4�e*'R�`�3Vs�#ą��|w�g1����ԫ��rB~�:��B���&g�c�?��'�z�s������OB����ru��,g�O~�V��3�c��+������9N1W�0Z��{��.%i�䘶|���Q�����1�9���Y�/ȦD��K
��N��6&�ګ�%�f9x(����F�+[���q+��Df�OoFr� �h�n�&�� "�@57u<�I
�Pu�*���2�3��Wd�}v��&�٣���&=�K)b{W��m��L��]/{��ܻ�U3{�B� �+	�j,�ۚ�=�C�;���9� X�0��!A�Au�+-����ɑ�4���e�#�Q�sra��d�����C&�%�Ti���o�v���x��?���	�c;r��2�����jc��������~�g!����Uj�ٔ:�>�Vѥ�[�ƲN���t����q�`�����,�A�z.8#�"�D
Xc��Rh������0�Nr:d���1Y�o�P������(�}�#X�5)�z+5TZ�e�s��
��N�+p�r�H͏(5�PV$SС���=Q��K	Hq�>�%F3>��2�������e��~c�T���w4=�J.J��<�R8��[bF ��Z��řE�-�N��K%��	&������ǥ7���<v("5�g�E0	��d��pҲWb��M���"����a���c:Tpq�~~�N��5"��y���Д��Z�Vڱ&fN8�C{΀�#��ʵܧ�Lg:st��yZ���̦J�e)���������u X��D�K3Xt-\u��V.	���/��菾�گ1�She �g������O�^������*Rh�4��_�ť�co3���������]��wĤ��\�c�U���t�]��t9�V���3�߶����'P��ߗ���V������Ƽ�e�� ���!0�g�(�M�������iSi�[F�X��Q���0��6p��{�����q(��i~~��ڪ�iOJ.����_�	�L��O��CW
!��d��g�%�:���;�������?�K������Tj	@�_�6Gc���;֪��[N�=��?��xM���lo	_b._���$�'�R�\3wr�����{��%5�mL�f����)S�>�[�SO��S����=zh���h��Q��C����G�ρ���7X�-!��Sl�q5��2ܤ����W�]��Y>U��&��@����e`�w��T}���K�۩�_�<S��.�<����P�v�t�_H�8>M�Be�����2OSRq�`�����+lLHL�Z�F2��������J��1l$#m"bĭ�EF΄9��a�����z�u�Ͼ�53�h����ur���Ţ-|�+L��D��;���C�}�;��	z����>H��="wrׁf��������wJbYW�Cߪ�1��pGұ��}0o$k��26�g��7�0H��7 �����P���O�xP�e6ْc��t�PA9��U�,�s�Ug�d�N�)0�|8�4(��F4�Q�'�k���Z��A�ty�0�d��H�r�˂����2Em��[U R����n�@u���:�f�ָ�{����,` �Z�.�-���c��� ����ԭ������b��������+X��{���U������N�v[Eɡ�Q�g��!�-��@��Dv\d%ٺ{�#~��A���-�Si���u������W?9B���Ϋ����`"6�ΰf� ����A {�����/(Z��e2J|{���� k��!�s@Ga_؎�(�������=��V�蝿Q�!����n��Á���Ed�s�]0����?�T�� gQ�
�#���y�������&fVD�R/�����|�H����Y}�6eOu���+��/�(+~������2�n�@�dt��#:��lۉ~�x�:�g�<�Cծ������DiUw��^�nCy����=af�$�
�3���V�=x\ifº�XN���2�U�	���2X@^z�]BD������j5��}+)ٻ�8e�f�tV��;�U3�IWL!
̚0&���ɮ�Þ��~8�Lx8�β�,�]�@�w4-��C��j�4m��������՜��Js��B.����L�2�����ߋ%\�ls$DX���f�[�9Rr�ݾ�z�����CD�N��
�����LlW�e��Y~}�����Ĩ��n�ʶ�˸�iP#�&e��
4Bi���`��b�Q|g�bq��|�I��1`%��`����-~c̆;�bO��4gP~Q�R�۰&Բ	t���
��jr-
ji��D�)�h���$Ha��ns{(ߊ��z�V��
/�R�t�e.9���h�	��L��/�,ȋ�b
������ǯ8��8kw��)��߫6g�#u㪭t��<�0 �y���(���p�4�͆�:��z�8����J�ι9�PS��ռ��҇}�y���Kt�
�6�R|��W�oJ�����ȹ>���wP�o&O5/R���[�2$w�� �g�Χ���5	��pz"��_ѩ��X�N��!V��2��/xdF��s4 ���//�?�
� YV�I�x��_UVUE��-1, �����R�}�A�"F�BAg'���7ğ��Q�]��ҙ��Z�$�ٿp���s%%�!B~m��\}2mቘ��P�91���#���2=MKM��r ����#��n���$�i�(���� ������p��YWNͅ���Q�i0�� �"��K0���r�dm��&�cq،rk+�Ey�;�� (�Ze؆��pj*,b��QX=��)� �֞��J���αRM
��_'��}�F����E����/X��y�C�@L*/�\ԋ�����Hϳ�e�fJ�������P��pC��G�5|�����/RDM��$��!�MVo�BZBy..=�G����<�����u�>���ߏM5t���
�\�_\آy�/cm<B�����̚1�#V#7����2���E���ULf��w�%W� 4�)�Uw~��Zj�7o5}�����u�eH@L�P�UP�`��U�&���y���e�Y�w*Nl�C�ԃ�:Y1���j�յ�� 1���Й��-N�������;ڣ�#GB��IQ;V�α�jF�a��cp@gvj�Ld�J��6��Z��K#/��ՖD��<L/����#���d��VF@nE��ǜ\Z�X<swT\ ��a� Biry�,TߍO�qD��#��]9�zMiY&�iD'��5b��i�>*��쀥8���E2��T�j��1���j��O�L�����u���#4x��A䆟�T��	��r�.U"w��X�+� pdz���Yÿ���=1˘I��N�1h���F�;I�ׅ��	��{��n���N~��򶑖��őn���X���r��^��(|=���ugfs����ht��w��WB��;
��cx�B��|-��2"�x�k�+|.Ҝ��@Wj�.�'x�Sn.!'MJ�����h%���I��H��X��a�[ �V�
��1�$&��\8�Fڃ�R&�d��`����B�P����љB4Q"`d���j��\u����O�;�6觉hM�,��G^�Z-��8�^���M�9o�&qR#w�2$�	��H;s��T�²+�M�Ve�`~��6�j���5��4'��zP�Dx2�d+��d5R�s7��/Za�C���g� k\:JNP3�Ϙ���5iV�(F)�&��mQ���[�hX4l*�$_�q�C���G$"l��<1_�y�[ �
;���Ͷa<��SM��=��a��Qc՛��%،֪�1�t=C��m���?�~�ۤ���c�ǽ�Xߊ�t� \6���}�[]�H���]��Ϊ2���bs��#����n@O>��<���
`ؾ�]�3�Tmv<����
>�m��J��$v�]ޘ�w�!S�c�I4֞h �̚����6)�dM�EGvC�i����̉�c�>�����|J�6�$.�u�x��ø��_;�<������L�~��'i��HI� -wC� �?,Ѯnu:�E��B/����jIt��t�] k�� �B��%�ZU��_��	4�x����ł�J�V>s.�L')iʎ�/��`9�AQ�]��%��t`.7�u�6�E�
��߾���fp�w�%�n9�\�6���Zx%
��X�i�Bإ�\_������ݯ<�
�K(��?�4��f�}Ey)��	h��)2�\أ�8I���YT�����y	;���D!l��cጟ�����N���0Q5(`�=�hv��L�pk^�Z�ma�M��f=K������ѹuo���t�YXK#��ػV�����G�'v8S� %�j:H�s���)�8p�}�$�����xL��~{����J$b�΃��%Vx�t0*�{������/�F����14RI;Ul�:�I۟�rv��A��Gv�	������M�v�(�>�:^�ib5_�6��7n���:֎t��W�I�p�"���5<\ [����3�%�%�:�����+㖋
Ķ))R @8"Y	�e�l��fl�_0D��>[���m������C��Y�$ʘ���>T"bM�"@|"��A&�uc�pd��zV�,�����iN���MK�7M��v��IeJ��r�F�,{|�x}�)�n=��ᨩ������M����7������x�q��s��GKJi��������uk���\IS�����t�wR{�z�� 
�G�Dz�o8�d���3�G��s`k�\$-�oZ,�b.d8n���6O>��w�Te����t/��َ!�7�_H4e���?��$K��4+�&�^`:A^=�#����fY��R�-%�)�
�}�]wWM��y���uᦔz��͓Ĳ�2*I120�|��c�I��S,�	��FE��4WVK��C�7���h���4!��`Ͱ��;�$\�nu�to7i���g�\	��-�_�U���(^�b9$��f9N*������ڕ4�Cܡ�}�Q��P�P���S�O�)�p����1!��X�9-���O8T�*�#5j�Ә��c+�c�h�E����*z�1M�UgD�n���~/d���O�{�D�*��g�'��?��B�?�W�����(t��l"�(�'KB��݇���ȿh_���D|��k3�J����N�{!����L�������t��M�rm�*U��F=�K*z��v�)ˆMX�.Dyoy�b�[f�� )�n�Z@4��ǽn��1�0�Sb+�:���VS�R�2�ȦGA�c�I86�$bea�N���Z�ZI(�?<��To[�;u{6ë}u�n��B)���^GB�@GO����W�+T��R�����?�l?OB����	�zJ۫А޺�s�'��:�ԇEX�hO��8:��׵�-�NfaƎ��%p8�E��d�ߊ�C�>3 �x�24�y�/��ϐ�/�f?y�3l0\,������6��*�pV?/n1���kX�CU��ϱH\�@W[�X��J�;�ba��ۄLy��� �Cm�����TK�j����bA��T؉��v6T06=-�:���4`�k=��G�:I$�9H��?�O����e$PE��+녖�iD�e�<\	�U���9;�$�2�)��f;�d�9��F��k4N]��y�k��Lz���7��tp��A4%jlvaau��Õ�P��>���q�t�����K��P��fnG�[p�����#<9�8�D�c�NRS����ÉJ��x��J�-n?X�c~;�Q�-����e�?��!\|%���"��`�JZ@�h�#���Q������?��*.�r�����[�H}V��xqNb�Z�	 6��T\�X��9c]	���z�=i�K��Uբw��;�܄>���/1�Jpx�Pߑ4���N�����_�M�t�<4�9�(K� ���%.�a6������7�W�V�q��76��鑝;2���k�������Ph��
I�G�Y�G�ht���*����<��y��ؒڐA�N<��ʁ��1��+�OԤ���q�<z�xD�K��N���t>[*�؆���=�x�B�N��$3vln�4�c�R;�Tv[��[#"�v�q#a�_? �Q9�iRP�����YY�� "�<Z��Z����T���_�~X$�!C8}���>����^͙<����bs �VΉK�O����s��wv�\bl���.J�E9�MGH�̺ �d�|ID�`]*�)�-,u�����/�����p�pK�ޕs����&u��mU5[[m��2� ;�H�ߌ'��=�u�� �{�Q��N��e�������o]��܃���O�%��~�� �m-*�@P��4L~�"���p�DC�#�bk���7��t�u�w���a�n�������_J�ÿ��ۡ(j<O4�I�m)O��?Q��AA"H���Yn$6/���a�	K� �xh+1��r�^�}�t�à���Q�~�쿶(���7���'`�·վx
�����?��T]&��]&��sS�}y�$<���`v��v��A:u�	�Ҹ+FΧD�~#��@�	��Cxr��$���In��&����vAچ��W[�Ln �����ȵv*�PS��TV *�Av��_S�G	�E�_-v�Ǽzv���ڷR�ծ�T���)
�n��b'�������V��;�#إ�cSplJ4m��Rۀ�h
���5X�:�'���X�ȑ���!-k�+,%��߱�:�q��!\"��Hv�x�4��{T^c��4�t�IMȆ������-���1dY�����z>j͙�uW���T�R(M�DZ"A�Ʊ_�@����[��W����?��KQ� ���v�m/���>�_�
)%>~Z=��P=��)~���d*s��X���ߣN�y:��bf:�N��6��\�vI;���q���e�$E�>8���C�Y�i�{i��?�`f�ީ}����g�d`�E4e�/�x�޹�h(�ȅf��h��G�2�����.��%n�:�j{xӼ����w ���̣�ƭ��U��v�)�|^��2۬;��v��L���S{��Q��)ˁ�_�l���c�Q�<P��+0zKO����S�#Q��򍺾V��f6kL�`$�a�S�:+z�p�y� Q�g��q�>z(31�Z�/T�R����!�A5BjHǚ{ׂ���0�|��Dc�:��)L�p���sc�c'8F�U�����IZN	y���J�k/gr[�,^��K�|%��)[����i�]3���X!�{��5��
v9x�ĵާ�n�V�d�bK7����9�-�xZg0qy%]�&�ӡi$�-`״J�d<1\�O+��dE4�D
�F`1������<��7Ҕ�Դw'����dB��\9V��!/��V��]f�}��#j�дzx�17w*�������Xү��.�ö�}������.2S�4]f^v���v�w���B�P�xY��X���yrz0��d���ʘ
\��0�-�������;�%�y�ĽE�����0��&�>pߜ堩�Nl8�Y��)+��|;���q�c���֥9�j"�Ӡ)�#e�A�έ|Ԛ�w��n��7��e�L@����%�]y=EL�ȹ͹�&��*�W��*��Q{߱h$�mӸ��Ű����ё ��u�K����+�Bť�p	�$��b�Ú �ua�qh��\JaF�;��ʠ&�uD@��%I�=yX ��Ӻpi���g��1S �{��hۉ�<�^S1j2�Y(G�~���-rs9w�B���v �C�v�4�Ƙ]G���B�!V �M�X�4�����{�8'�zO�&��zﲾO.���9����Z�ޓ��%Z�F������uq�=g9b
�x���ixD%B-�c��;3<L�P��z"��9�s�����>��ҧ�5��E���6�˗?����)1zp�5|\�%zD)��;>%gR<�����Y?�33��6zH�o�$�����s�;�D_����s�DY�?�>� LE�
Q/@��V�.�T-��E��<jv���-S`�Uh�h?���7�N��n���q�;����æif=�R5q7���V��@b8ԞC�SR���P�WKG�U��:�;Z�� \=f���bkܝ�������M� �+��NN4��g��ũy��hN`��&U�΢H}�٧�DʽY}m#��.����09�Jq�1#�^�Dd$!?<~�maL��� 	zB�7q����Hf��oF�3.��$JZ������Gr�
�$D��p�&���0:�[����"��1��%_ʣ�o�V���y���"��+� dX�n��2� �X��W��Ր� ��3���>���|�,Z6�-r B_��	��I!ߏ��X)��u5�Vk�-���\}��ˡcV���U ebB�����TQh�}�}�־�!����\��ʧ���taU�kn�bH����lZ�^`T�x�� ��ި�d�ʎ�'�ޥg#��;C���c�ܖ9��7���dRm8­0��du�?����E��b�x��K!�z�)��<�K��4�:��R۱)1���p0��t��Q��B���5�?nX�	9>aVT�2����zЂ��~f+�a�Yo��+�������B# -��9�DÇ�v���0�s�$��!����@/ˁN�S���ؿ|�A�hK�Q#��4Y��hSR�MT:����M�q����j�%Y�s0e�����P(���ui���h�$ �u�҆�=��w$HS���H���\U�l�[|.�����1��r���B�)`]��U��ݯ�vF�g�m��}de��t�%���
S�������&��R��6�Ol1} z�����Ec�<��0DXʊt�%�5ǫAv��*3��odظ�M6TB�1.*M9���ϲܚ�C}�8�Y��7�_œ͹�IJ�� +�lb��6�D��ቹ�������;�Z{���sP=Q��bS3�GdP_�x��k�f���*PC�z⇖S�s4��߹��*7(/=əw~�By��> 6��Y�"���@�ր�ݞp��/�ѳ�+���F���4�i�W�:�C9���r7�}��H�>�f��8{��� ��@��䨊%xs�"�c�?�\'�<��v
kZ�x7z�ul�V���h_P=�=d������4U�9x۹4��3UzCxv�daf�F.v�����NS�Tz�+���Hc�n���������g�����čhA7�/��c�;T���Қ~I)���ui���6�G{�(���Yd����qؘ�����N�+���o{<�)9��w�x��*R���O.a�&@�En釰��-�:�B�(�e�M��w̓N�i�z����,��
��0vV�L�ihxtO��=+�0 K�TW��� f�gl�D���g9���fe;��&���WA>�;}��a�j�c��g�Á[�:�����յ��O�Z�(�{�ҶR��A�����GŜ;�/�S�Q,��{L�G�z����҈�yEx�6�'%��Fr:$�bum�0Dk�Pf��4Vݬķ+�5�F#{XO_����������-A�_{ej kK,=9���y
�0�+����,�r��{�$��y묖}�����s���F��ƹB8p��_�G�}��i�������7T�VxE>\m�������۹�C<���Yȗ��B|�᚟Ѥ#3�NA8�m�7��N��T2����j�	�f�#�H��n(�CZ~s*�Od�[���?�i�:��)��H��R������ċ:�5�Gq�y2�.>��HĜM���0-N��v�W���ˤ�M�quz�ˤ��(7�S�Q�?�%��v��%���߽6
�Y���K8y�����|��|83w�P�O�e�"||��t��*[N*ޯ���	8T1EZ)�}��=�����HfW��v����mgg�WY7�\@V-_��&}F(���G��8U����/��AU���cn�A���b���g�6�x��>�X=�����/�x��ZW6��;�f,��K,>�'@�_Nڋ)7V�5��0�$�&	ӫ�ۯ��C�����u3b�������{�X.���y���S�?quϋZ�,4�.="+!}�dw-	E6��D��,�ek�#[ŎF����k���X*Y��)��̭Z����=5��6����	K�R%F����g�i`��l^�%xn4�F�{(�E�H��, �1�<֫�����z�oD#��[��d���yɬ�Af�Vwy� ,����6u�X�3���n�N"���/�2��@^K���9z��Y~
�,R����D>bF5��ʨ$͢�#tJ�g�zKb�?��(��߄MP3W�q����G�$${����|X����`��ܾ5c��cc�j{��L�,%���)'��
d�_�$M��0`l�O�^ S��<�~l?��I����Lw����b'[T����ܕFa5R�D_.�k��|gK�깊��LD�}�?���E� .�|_�M��ɛZ�� G�l$��C�$�!J0y�9@�;b�a )���#�Y�-tL���$SO	8�?�e�/$�]MF�w����2�Ǘߎk�~�!
4�"Q��?¡���jI4�ȧwjd�/h��pz�o���o,lx��H�2I����x��ΊM�'A���0�Ԧg�e| �޷P`��5��}��R�2�J�b�����l��/�e�b�6��Ў�(�)c��P�*�[�7�X�&�1="��ر{��P�$&Kz5�)T��~r�nK���W���k6r�zV^�����-BbC`?K� &�#sV���v�˭qQ��{JdPvZ�h~HOK8T�V����5U��;޴�ʹn���kRJ�WW���x��Z�9/*�z�az��Q� V�7��L�C�F�S1��[������t�AO�A�.�Jvɽ1&���q<�:
[�5"��Ö�#HIM@<f)�VI8ۑu��2�����,�[��v�*)��Y�/��KO����S[�c3q�4�t�ǣ�e����:�ۄQ��
��$�s�8�z]f���l#�j��/�X�J������8���>��?Ɋe�
.�pvb*u��ԭ��q��L��ȃCE˲�Fr-�|���gw�c(�qƮY��+H<:3��^"���������CW��SQ�{trOu��$�n�P���
�0"�A��3O�a+Xcv��<�����Q�8���/�/3@��Hc`���� �-�7�碍�(bF"��l�`l���(6��w+;�^VG�ߢ�.U�)��e;߬��;òS/i0���Ep�e��Ӻ��,kC���s�z!�[<���4ҭԔ�m�YQ;��3�xŕ��~ߥ�ue��.}d��0��QL*[��Hc����ώ�s&L+������H-?v��C�u�癟O����M���O=�T_���Y����� 6�В���Q'.�Ŷ�!�E .���ugԣ� �㝧T����$�^|�WrX�Pn0�CE��c�
!+�&Y|�C��Z�R�D>o�&��
w�Wz��;y�_ a^��b�5��P�;.�&�m�W����c���h�d�3	���v�}�yi|m�Y��%��4�<��vԷ+xo�CN�G���c	 n��G!ƫ8���]|��������m=z�A��M�NP�=��/�U��!�a������\��6T8�->��X�ARy� @�I���/&�G�?�Ҝ�kR����u�� �d�@�u��uK��F|��PS��Xw�b���	6�-� �]����y�����B3�!3,��]���~[��;SV�B���9�B(��WG;�ïu�C!-}1䖤|pgSP�H��^h��M<bp��e*�ş��j�� ��¡M� �*JKT�����X��A�s.D��>8���M���G�0vc�P|�����(�`#����[�5��t�Ͷ�����(�Չt~G��9@��9���Z(G���2<>�U���/t�,�r�&V���ceb�)����<j��쐈�~�&T�]�Fgo�.��LS��02�n6�^�v�����z�[�	�#����<�lߏѢޞ�����Ƣ���($GF�m��Q�{�-u����w�KHl��8�t4����0Si��{���z2�d�+�+L����
�a?�-N~-f!�fB^@&��;��|jx
W��U/��X����V=��-���g;�ኵTPy7C߃���#��z�������W�(I� ��3�5�ό� ]3tR�e-�ܠ��-��k>�٧	��"�p�z�@�Ŕ(�l���7@n-�������Z� ����Bonbb`~>�X���[X�t[Fv2��X�.%a7�!�'��ֺC����RΧ؞�Q&1?N������]-�p�/=?3Y�1�H$��m6�V{-y9ܝ�eu^�;ڋ�w�;M-�0�}yh?R6D���#p-z�P��XO=�4g�)�������jf=�`v����X����)���L���V�`��/�CN6�t����2�v���A�G�	V6�k�:k��T�){�Q;¤�=���3��M�Z\t�1y�:`��zn�u�bN�&R�d�n>i��}�����qt,��q^��6�~e�N�m��P��&W'k��7�-�:s[zx��@jyY����T�b�Wb��uR�� ��շ%(�`)#ṫ��7���y����m����~���"3#�R���˴[�*�k,��m�f�̽[Z��:��~�I�-w-�fD[4Z��k�?�hƵt���|c��	g׊d,�Me�Y�^T��1�!�G���_�	�B���|��s���#�O��2M�e��������u�O��q�@���v��O����/v��a�y�񬕓G�1x���L�>1V�_�Nd�@���4�h33������D�Īsy��UG�c�)�����!YN˺����2���u|�Z�q����zԻ��ƫP��[Xgݖm�,L��el��CA���)�뭌~����~��u�lʅ`w��U��۟
gBl��ll��H��/Kh{Y�l�� ta5�x��Fd��噠T�Ћ�&=c�Z�)�9���Q�X��c^�su[��E�=��Q"�� t葐�0qS���P|�sL\c�ޣ+&�)�;-�gWXnx�(�zoD��~�{ǅ���8��`�� bYNu֢/X)�Ӏ7h%;�怤X�B��u�?%2�K?�Y� f"�U�5�/3�P�m��ez9�r .�(c�0���s*ڔ2ŝ�D?tM!y]F#�:���l��+(�D.MR1�&��$�S/eiY��!P&3����dI7 ���mk	2����ÙG��C1��72kU����<\�%�0V��e�ؒ\߸s�T�X���Z�Q]>��-E
��<��N����eH?$U�S-��$�ec��Kl�i�3��:������zG&��C��= �/ɥ� Q���0��O�≅D��Bq��Ϳ�ش�*�\�Z�������I���L�3�[J&���ݟ��*�v4���#ٕ�+1�.>�ج�p��,w��kvޢ/�U2���^vi�K5��b(��sQ����)�#�Z�m����~yZBK���ٮ���	�#xâ1"���J����v�����rܥ�aq2n:TiN�~��o���ڽ�k(����������H��d��[G��=��wK�gب�@�:I���F��4Cd��tu�"w�!�����M�Q�G�L5VFlxb8
AWݯ�*yZ����^�'���QZb��	ב"f�������`�RbO����%�宍��O��|J����}���D ���X%���k�T���:[G�g�~������w�\]3IQ�F_�]&L�N�g���t��������V�u��US�z�d��M������/*��&7�m�w}Lk������2�`v��d�s�rûp"�[ݝ��MI�?~s���U�/��ޛ����t��X����ټ�����m�[���:����"Y�
�(����]����(��B5u�����$�z��+��q��u��у�KV�j6���|2�wd�����J��`���w��"���iH&�WH�QSc��o|�� w�Xxl�k�qr�ƂV1Z�.X�ډ�Xf���f�d�"20b�e`	 ��}������q�W�v	j��iGF�(�τ��x�*D'�ӛ�� ��Z��q%-2E1�uݎ��d�� �$�2�p��]��g�d�%�Y��u��ߚ�����Y:Q��X@�5�]�'D��x�j\~ tX��7��9@Q�8����0�l-�Zߟ������ԡ���ֻә}|��ů��A^�j���,x�\���Խ�B���9���S��>��l� B+�4���D��)yn�sӒe����s�-������6�n�0
t���S�����=V*�hЌ�i��ʂ���YFB��o@KaׄD�F����aX5G�i�?�뛖:$�<��J�?�CKc.]B�ԛ�Y��p�!�����$)�\I�SD�7�0�7�);M*ھ�`s�)e��6��h��uZ���(V�W�u�#��c�VV.bk����i��PY�\ z)����;Bj䂁�m�s��	W�[90���$EeXp+Gu���ռ#-˨Ѥ�:K��3�Z�I^�bhf�'z��?u�)w�.%�ʬ�N�=Kp���L��x2��j/d�P��g�?6hB�����i�nS��Te�^Rx9���@ Z1�7`�
�� �Z��	j~��U���2>1ѽ+��R����>��06���Hэ�N��7)�������+|�7��Q��~���0A�^�, Z��ъ�rzu��=pZM�(�1�f���ҧ����G��u�_�ʾ����o��)S�� ��,�n���n?�MA��¨�}Li���,������b�R	�1뵿�@7|���1h�`~�'����9�~��C9w���W��t�v�ȷ�#e@���0���$=pd~��2i���-Y��
=/����.��R��+�^�'�F�>�녇�9kQ�1�mMɾ[4�~{̸D��8���,�{>7�Ԥ�5���U�R�9D(�X ����N�q8,�A�r�;�^7ʖI�Y��_5�o�nt����"�K��P�).����6�p��&������ ��Bu6��Q�!��?@A�p��Ƶ	����� �v�>3c�]�N�����PR�u<%d��]�u�`k����6 T�}���{B���P�'���ƴ�=#r#'�n.�0&�.��������|V�1�.�;-m���LL7L����O���\I�<Ԋ{�Y�V�%��,He�K2V��X4��>ĝ;ӂ�z�
dFǁ�i�j�},s���^�����ՊvT�'=�2�xE��po��ju�6�hEGh��<h*`�-����7�<����_����z�olj����p����xm
������7m�k7���X�H�t����mI��	��l6���tG���An���&<�#x�R�2g�7�ߩǻ�9!��QW*O��J[�v�}�k�۱t]���Q��%�	\���j`'V�y	��/�2�u���X�����#��.�K���*Y��9�Gǈm}�&gu\¿Ǒ���ɑU��%�<�r���ϮeS/��_�OE��a|%�8剏-X�����mQ[��q���_��0$bUT��N�0}��Wc U�șO�?�4�ؾ��K�9E�۴4'��}IG	��w��0�)�c,��8��U"�)�u%M��⯃\�Nq�����y�6/���,����
��bac�� j>�_�#����X���t±	�ɵ�<��aJ�/�>p�u�8Q���s���μ^�3۽j:��������ۿ� �P^֞b����_K�7�|���n��T��<��q}]�&���/ba&�b/lY��)�����LT�+Ƙ�i�/��o� }F~5]� ���o�0GYB$����V����s�h���
#'��x��'D�0��3�*+4RD|G%�X/�8�G ٮwof�(al�﹊�C<r�7��e��xv�~%\���_A&��^�+~���}6�_�gR#��}�FwA��MI`=�#/���Sɀ�߼e E�sE����c�R���;�S�Ԩ�q�B/�U ��� ^"�bb�V����+51�«-��=���4�������0*!������g
D�X\јI�k:KC{P�h�/E;�Bt =p;m ��-�a{�l�W'�x�;�ӑG:G�{aȎ���TW��}䏡ZY�.���8��g\_��l?�����[�T��0�[(���6s�����5t���m�Ke�s�����&JYw"M����oL�@�l�["T8r����|�4���	�=�-ڛ��6�'�l��[�*w����:�[�S�l�4+u����}lsj �>�Ǿ?�8�]O�?Ά����`\<m#K T�}F}>���# P��[��|��[?̒%ȍ\�a��9u�vkp���+�Smѷ�[S���,ev٪+^9HO׮��y����:)F�.;&.!�Ui��F��
�-�.;�omSҫ3⧱��hv�p����OF�����
����d�l��̈b�4�*��_�!Gy��{�α2nIM�w[��u���p��#�����=�,�{՚$����9<V�ͮ��H{T���a�a-Փ�$
YSӽ�~{ �O�Կ���~+���I#^�L3k����/��ۃ�#��W'�F�~�N��˂��i j�OW�᎖����2��T�8�8��A��da��r�1�nm�:."���Lf��'�"	G����O�G�;� �5�Q��g��M�2�[d<w��"mȅ3H5���22����=�c��K��Y�v�a�w���T�둓]�����!�����b൨�|`*<�@��5Rt��c;=�3�ì�s�R�o���.uU����c����(�XG� *sXR�	�'xJ�t2 O-�E�v��"�B������{X�8&&^�y$v(쏻����%��ٹ��E�;�����_qt��9��`�6o�3d�w{�][�����X04<G��^�w��^�2�G~QA���E\����/�t20^0?~D��A2�5aM�m\ea$� ׇ$B��_��v�44j/*�9��Q�t���t�CSp:�~:����o.}Od��p�[-]0�S4r`�q�������~cGEc���+����hy�y��R��.�s�FQg���z���l�Q���� �r����k�n������f�5h�v���T��`���Z���s��t/V/���M�qܞݳ��dӃ��Q���5T���n�
��s�RF����������n�ܶB�;8���ƆJ�T�.I�Y!#���CΖ��Ɵ���{��F|�`��db�O�����/�8p<+}Z��O���Jv�@=ur�3f��"���q�|`����j��	������'@��y�}��	�3Δt���b�����qUc��gĲ%P��g�H;�����Rh`���o1b3=F""Ŧ�y Nfp�"u�7.���&����"r������@�ׄ�SLC�"�3ǐ�>���SHzb�6V1d���aF��)�Ҵ��Q��&���b�?Ըi�xh��*'`�Q���o��@E$�嚄�I�I�?��}Js<�6��ʴa	Ü��rwvT%U!��"����� .=E��C̣��3��HY F��1!I�2��Y8��Qk�i8x�� �.iH���,��k��-�y���L�@�])��B\�i��uQ��W������f�'7�l4ڏ�H5b���f�,[��+�L�k�?��i_��z��2[�e{�s�ǻ�=���I�Ƹ1�n�	�=?���G��3�S�B�C�������M��N�Y�e� v���[F{ޱ[�
��Jyp��1�\�9</`t���1*�/��@�YQ�t��df������^���s�We�����9 ����ڤ�BN@Lθ!��@Pd�~Eo����f�\��qנśY�����5����:�`�E��_!�74��'�ә5�{��$(ܚ[���͸�>�W�������O�a��o�]d��Eـ3�x���| ��ϟ
,�%�~��H�\9���2'Sei�$�un]�Y�b�V�eO�ٱ¡�=�S��Y"���pUZS�g�V�Ά��Γ��M��;����%��
��\ײ�s���Z�e���!c��V��srR�ϥ��ԉ���J��Qɳ,Ս����!�:��h�o6,pMH~��(g�{+lK�N�I��ܖ��ή�B��t���Ě���]�����U!�z3�i�:*6�[z<�V^�L��v����^��T���2�5�Y.\�	������p���M�};��K����Fy���'\ӕQ��^ը
vk�XA)O��,pГ��v2��\@ĸ��Đv��w:�4�����lO���+ �������3����I:��n�
=�4��Ϧ��3j�4V��z}��esM:��#���o&ŗ�]������62Ε��$$�����I����F(�e�t�:0�r��*�N:jP��T����u~m?ц��s��œ���sQ���C�1�ʠfa�i!�" $ڍ�l��G������Y�Wϱ�ou�4�D	�}�=T9�%[mt�!M(E�~y��]�R���Xb�!�{���=��r������O׆�tjRu4����U'D�-��t��F �)�7�+���^�hi�aR�[��r�tݨ�b<����b5ܿp����x|B��2�bf�����>zR&I)��b;��%��c7	�|1�	�t�e	��қ4���vw�t���T:bX��� �vº79_b�,�ۨ���
{�D�Iz��;���j�~�6Ԁ����W<TreƸR#y����s�ǯ�I�lG��Sr���H��˹�B��M\D�+�8X��>�e�H��@�{�5�q���O�x#r��K����X�=Ł!,öe��g�Bf����)��e�;0��������xV4i��w��ڋd��RfwRc	_f'EPe]�걯�\%��3	ܫPL���v�X�\*�{>�~"2ن/���1t���WwgY!@����X��ҩ`.�ND"pH`J��b�]��s�n	�s�ݵΘ����dp��6f�J��9@!m1��KD���jZ�Q 3|�s��"s,�.����@_�Z�1�d�"��VȪd@�t�u9���Z+>���)M��?;T�N���蔞@I ���)O�' P�u�Z\� I�'�Ѥ����e��
|�^������	�vh�Q׬�f�MpHU6�� �tt`'����`�+��H'|6�g���&>�k��0�9E٤t�H(�6s���@�R�E�m�KDd�yđ���Σ��u�%3
�]��O���c�������k�g��0���ڌ���~����2�r÷#���P�_`�)#����<-x���mQ��Y�=h5n�vP�"w_l% �;}Aײ�苃o�ܞK?����ҩ�MC:QiB0�&.oF���8N�0�s��10^��qUw^p�XA-pv�,4�ap6�Q��-Dg �(�b���m6-�}�%}1�]�L�:�\k�gJ4!w]��W��n�|4�Qd�	�
��)��72P�+Q���'eN2�^&G��cYo&�&rE���ϧ]E����`�Zo�e�;�?l@"Ԑ����>�E���%��w����R:�4�{�<۷���~�kK�={2�����A?��7��I)�KR�8Q~�$&Gs�_��W+I=&J�S��Fv[ ='˵Q�E� �.9%Q�U�Ԩ{| 0s�j�73 S�f��3�Bs������ZV���|�AI|S�z_ӵ����dZqT��#6��q���bZ#jP�J׀�����;,��R*�,:���Z��,l��H��DYP������J$�O�D=י[�Z�M� �0�3���D�V֝�	�,�{bs�Q���:��=Y'Rw�|�� zS�X�	�yExx�1BW�hO��ɂ��_2���K���9]w�=N����'�1��q��B8�/�T���!�J�u��J��-:��ۈ�#vF��c	�ӣd��`�8T���u�K_�/��x�l���gvj��Ѕ	go�gS�{���Z�#�$�9��4 ��T0�[�9kT�/lw�*=��[@�j����pw��LN���÷B�5 ?e/f	�ĦZ.�w��3��F���'�]��[�"f.���R��KY���{�~PL�j3�3F�1x\�����&�qt��$�Y�٢ȃqr�|6�JOU��K�6�84�!h����4T�ؙ��P��TQ���RD[�2 ��{��Ѻk��׏Z&�K��Ѩyj�l���|������o~��Z�	�ҕ/��c�7��c|w��RX��W"\�J��c��{Tc�t{%{]�*s�������#�M3�U�1�u4	�*���1����(D���|�I��mw1��
b;7�K���J?S�!f��Nw~xzu�#!��e1�WX�$`������F���f�S?fP!c�4E�!�,e��׷-J���d&8�7�����gl����s�䌮��<F�g��-���p7^	#W�uu�^��#�۫[Фt��ZY�9#��;�f˰�3.M~/�\$5�≂5
T0z^��o���$<��Cww����A\AX�0�.�U�;�9~)qr�Y��!o��o��l�<9��?��s��V��/b�A����� t~�M�zX������7�w�����=N�_�O��l{��@�3��^f�0H��S8������:b����Nu£=f�`\\��#뱢��0��ݦ��Z��ZBr��E�p��嗶��������>Q�.�6�.�36��p�Ml�櫀v g��^B���B5��ӤT��u�.yMK`1�0�����g�Dr>��FRJ���������O�Ј���G歟�aI^O�
��ǻ���r���d�:���,�NMA�EI��׹��gdD[����2�sc�w����~g�b���m��1�UHG��J�Q��O�ƿfA��TX�j�eca���9��_�\O��E�V�&R�,=CJ�eI.�iIg�������Kt�	������5����E��\1�)x�h��(�V8B�r�=H�O�������y��1O����&����y��8�%?��`�é&l�R��5�!r2Д��6]o`Z�T
���"�-���I� j�CD����]Ȃ�ʸ:��E(F��J��9$i��z �T]XJ� r��VJ��c0$�إ�&Wr��iE���Q�g���f�=�@vG���I��� ������W,j�0�&dk�%�Es|�S�v�k�����1m$l��OZ9���?A�Y#�*�vi�E	�,�o���P��N��>���*w��e�ߟ�)0����#��r(}��.���&!ĵ�U�AlR�+x��q'���"�g�iu�z���UR;���d��B��1S�����-�b��88�=Z�3��t(��s�UZ�9e��m���=vO�U�]=�@���
{�'8��e$Z��$l@�&�Q��\������[E��rn�����H!���:��<_�mn�cNٌ(�Ifm�; �I�U2��n��������H/*� �8蠏g�1��^�B���q���܆���#i #L����7g����
��WX/��MD�9���1Rx=o��3�G�)uSϩ�[��y"�G�и>=;y�W�uջc,]7)f��̽v�hðA���9`) �������d� ��y�x��V�ҥl�$���*�3U��Y��k|K��^�Jdin<;	���B���}@~ێ����2|�w�_���d���v��L�3B��s��P葵�	wI�����@|�rf�5�֌��CVώݾ����"�~�aK|(�3D�ݾ��N�B������,�2rQ�v�:�5Җ����3q���b�~󗦒�J#7�ڜH�*�m��SHi��OXϔ����O2�5�����#�������ņ�:z���R��:���(���7������/CҎ����E(��Iz��`�>����(���B�6F�����n��������F�y���!z��;A���kH:�睺��<��U-���$~����<���"D�y�Ā.�՟JIA�B�,��]��C����f�l*TÑ�R�:�S��U��EL"����9�Q5o�Rf��ؐ�b�Ws>z�l��}024��[,�v�^T�c��Q\I>U�M��AkW^9�%�v �P�ee�.�;��u��?��c8��o�2~{b�1�t)Z�=�Ӯ�N�"�+����.V�%�㰣ʤ�-~��|H��WП�X�E�#�Ms�5��`u���@��XK�,���Gc/��̱T߄�S��:}�P�X�H�t�#T�gh��s�Cٓ�NF�}0H(n܍����Pe��H	�u�F{��s�\�0x�)�e~L���H)`�����Y�! �O�X�=-�x��i/*qwP���X�n<3:�W)�#�������H1_�����A��ac��Y�h�G��b)�'1"�!�dڿ���M�$	��^0�]�sC��@�:CCbP	��$��X���Op��KĀ�O�T���a���"򱻼�<@�^6{����J�vL��
��-l�QhS��^)9��Ņtm��Jk�<;;��,�M�4����{���^u�fl�f�}�ā�	ŬD5u��E�.p���
}�h��T���t{�-�9�~�t\΃��'^�}<�x��t��ar:�N�U��~b�f�&��P �I�Ռ��T���E6�4돜t:~��$:o��x�]�}Jqٮ:�mu ���k f����(�q~��׆���}�0�/S�`�+���2�!�i+]O�Q_�HR��m�N5�g3J�h��ʩ	�t�m�jT=jX�	
��i�]:�W1�bVg/b��=�$�rBע����LMe�+VE���^J���t��QdMy��q��!�.��P�E.����h�[я䠜c���hcuEI"�Y@�[��+�N�%�2L���2ha���������us>�J� G����N<"=.°)ɑY����C���r�u9j���b��d�t���~���{�>�b����a�ߺCA�Kb�ȧBD)���C����ˊ�c�\�����R���:�����M ,��[hն����'$}��/	A$�ku�4b{y��ȇ��G;�v7-�ܪ	"�C�q�����i`2��F�6��nW�Xkn�^&;&�V���@���¶��׈PH���Ŋy�'�9`r�0���u��^Ѓ�͔�f�D@��L�1�Ut����AK���8�1tރ��zi���:=7�5�tڇ��Ǝ��;��7�Ñq˭��"����q�7W�)9'�Gm��Y��� <����Dt[�Jܯ�Pg�QH�:�D��Q��u8Y�uȪ��LB6)8qyT�!j����:	P�z)�T��|�&u��58b�%G��y5xO��M|?$'�;}uN�a������8��5V݉�w���g������ �`�P��.��H��P�!�]�A���oTO��$
R^�4%�6߃Q�E�a�C�Uz���lo���	��&�XNf�&L �??~9K]��bJ������ۘ�;3ؕ#�*د���A��S!z��U��29�����ܯm�a��Ǿ\�䒽�bj�d�if�)�M6'3ϋ��t\�?\�O��Gn�a
��|q�;�-��u�L�f&��N�z��/� 
*���
;���4��#�K�D���ȏL���mZ Bp�@}pz��y�X�"����"�teL'�`�&rn��W�q`!�s���v���Lg�fG&Qa�o�"��u �<]��g���}�T.'\Li�i��ٛa��t��D���4�Ε�����l�c�rk��ӫ�|�Yi�o��瑔@|(.��(����C�<���ُK�Ō��q:/��Sl]IU`�#�2(c�!-?������o%���B�@G��J�I,�!�Ev��ȡq�⹥`������C�讃^[�h�o� vBDʹ�0�FӒh��cWٜ�j���w'Q��9�3�F����L��$/�5��Y|;��;��G�J�D�cҤܜ�w5! p&�~�-0���-R�et�� �h�z��2L8U����Ƭb�Zk��|Xe�g�Fw�A��[+En�v��9�7�%j!bNK��z{gZ�[ �vٛ��%<�e����;5����J�`�sʳjχ�;d%�R�9�a$�x}ߌut�4���T��²Xn��!�?|��q��ɖ���� o)Kv.��k�C�=��,4po���GA�Z?��C����,Ca�d��
��2Q��l�j�e�T��-�B�^�����G9*�a+�m�kBk<4��Z�$/6��#4
�V}��$w	���L�A/I�����ɟ"�3[!X��r�-I��`�-(�`��G�7A%�v(�V���rN%<�-;ª d��<��e�����)&V�K�����5�{�ˁDi�AW �K��`EX������>�ǲۂI��EY�}z8c�e��	�G ��P��}qSqD�+f�?����X����_Yp�Y4b��/�%��b3�<dX_}�ɾ��[�X�E�Hck�6b�	}����#d5��t����k7�j��ӈ]�^9��o�����I
H@9}�<�#�O��<�cD����m���?O����y��P�W�m�-�j�zn2?�9�G�ja�3�s����Ś,.�Qp�!t�r����K���_mI�P�I*��I�'}wͥY�zė��NY[=��G�Ȼ���F��Y����젴�=7�*'ο5|��){���ݮ�/Ά�S�'e�4`����1���9�uSW��P8%���ejߘ�/����t$�FE��;�e6W���l�|��D���-����g� �����_�76������H��Jlۍ����#��Ŏ��eFYϔ���,�����:�.d'�ձ�?�$(Q���/��ӇRz���0���Έߖ�,��}�-��ǽ %�eg	Z;j�P�(�j����l�2(/&��rTm�>��և�@}v����ķ���E�~�hd�̵ei&w�L=Ot%�@ɞm�]֬�*=�ĭ�(�s��e��V�jv����q�;����nt	���"f=���I���2���2L �l��!�e�UR���9�I9a��L��Q�p�(d~E���7��!6�ʘ�
����dEK$!6V�6�E�#�lQt����.���d[)`�|��LL!��?�H��EN�ƺP��M�L{��R��g�*r<h��d��@�p2!ʨ�g��~�Ty���͏��[�����T^N�D��F�̍��sj��+`��z����`�6�b������ߏ�L��3m�@�T��t ʢD�"d�*ͧ�a��\�rvl��<���ZVP��8��Ԑ-c74��mX����;4������M�>@�=$�ҏ�|�_��e$/�O���\G��Y����M��@�͌|��8=%\3x���<�+�2�=��h�U��^]3�E秩ňI3��v�w�6�@0��sD tΑ�T~w2�͛6P���!p'Ѽ�m����=.D��r�'ȏ�֛�GJd篿�)'�z߸JFYXK��p�M��7,A)	���8��
�L2Fb'V�DF�פ�����8zA�k9H��/��S|GW�[��1����<��Oe[�z�HNi����bKZ�i���"�C�Up��X��2?S��,�i%s=pu~�Pk��mJ�^/m�|��zDK��Ɣ{T��`�n���@1匠J�'�c�Ʀ��f@���`0���A-��0���\%d������ŘF����x=���Q�*���9ك�2��$�����O�����T�|��-��yt�o�~�D�1��!V��4�����S�� 8�-ќ܂d}QQ�wS/'�Fi��y���VI�J��O�E8��d;\�%j��!1�Vg���ūUݽm����-���];�Z�Fl2�0���"%�nb(�SV\È����=TW����Oǭ=�M:���m�+�-��~��8���w��ڡ�*����}%31���o�-R�j�n����r`o��Vĵ1���!���,���h˞���Fy�t)�)���j^�§*j{R���jv���r@L��Ÿ�y��u��9�uW�7�~�@SaQF��b�������W�q��6E��!�q��O��V���̌��(���e����D�A�Vp����
�|���if��֎f6�	"?�GI�9��
�6>���ă{E���({k-�� ��q��d�N0g�{iKzӶ��{���m��h�o�ޣ{�ͮ�FU�ǭ�"� T:�T�ӽU��/r� ��@(����a"��GQy��*#�}5�B�!�<��s��<����m��$l�3
���mN���?]��av��NB��"zC�.�e���^�����ю�us�=l,qg�5N�c�yM���Պ2�$癚�VO�H�#�	�o���sBחar(?��d��m��+h���KNH�����E5~�^#�Ir�*^�������3��o�w��1̴�4��\nS�'��+(�J�߇����ND��Q���U����wf�]5��Ns��6����3��|`�W���>Pr*q)y�����s���%=n��Mp?�IxO�t��R�l��B�#7�.�{���s�薪~c��b/qY&���[[G��iZ�:�e�:�"s��An�O���kiZc�4����f}����������*�+7�+�!����z.�Rk:��-w��@ �r
Ji�k��@�E��)�O�\y%rv���T���۟\�?=�
�à�`�lq�����o����1�T���e���z%uSj��XT���)h����� �a�W 4�>|� T�>3@uy�Cn�u�h奻��.�ڔv��vjJ�]|+�y�^Xl:Oe]�/���.F'qxO���5������USr�3aʸq���^9�!�-�tB�;/V��zf�F�Tڷ�����&=�-�l�bǢ���oy����C����ލX���,@刯���)^o+	
���N
g{������z/v�s��C������T��ٚ���8�$����Ƒ5��~2p���F�1+"���o�2QJ��દ��a�-#������Cn��&:��GVL����b;��ʠҜ���H�X�/�T��	9sh:ϯӪ�C<v�q�u�4�Kdwo����;��� 9i;��/��wW��Dsc���,ͻ��/f��޷��0{��^^;��V���S�k
���a�u�`ȗ��&4sq�!�/���I�]�)#�R��Iq�Y\� �YG$��Pr� �t�]XZ��:ڔ�pX���xirg���05����@wI�Ï���qb���L��Y��M�c�������W���&l@<Z��"j����%��i��2q5�-3KTF�36No��ֳ4��3������M{�O �hm�K_�g��a�I���}b|���a៓d�<���By�WcN֟��,5ե���Þ��Խ�x�D��;�Q��v푌ۇq����{�����+e��j�IFV�CS�^
��j��-���N!��*���J0���)|%�$}0��p��:=k,pجQ4�Ǔ!6�P�޹W,�m&�@0�pZ#:��<�h���$�] GU�Kߠ�%�yg���6a)�C$r��Z�Y5��"�=�k�����L�>��q����6h��6����sۭ5q��NB� �"�	�>j����e�/��4���S.w�%?R�� ��.����RF�{�ZXO�ݏ�z��K (���{*|���֚\m�6�T��4�B�D�PI���� "hCӆ������.ޑ@�V�����7A
�6캽1_�3y�4ܮ��+*P5�� �v���x�~��е�hY��љ����4��5�[�
��H������Dl������.�
a����������rǘ:!#c�W[;�~�� '?���19����@s�������C�m��#������ob�L^l)�@��$��X1ܤ�k͡4�)�y̟�P{� �(�C����''�A�oI���}�x,���7ik��K�7$�k���r����[m��xc��`'1�.(i���ã�}�>v�C�) Cba�i��8��`�G�x87�����������M�4_��~Ȱ���q+m�$�fh���@�`1ӊ���cfh�llg��1 <�`uς94�Ǫ0�=�1Z�ky��K�w�y���ŇYV+�����)
i�,��&��  2S�KԢ.BV������&�W�j�d�\:R��O~��:��-Z<�W�������J�	
']�&��(�/�0VZ*��l�篶Z�ig= �z�9+'�aZf��/���$����"����&�;xSp�Fjh-_���69C;zR�5��OZd��}-���1�qX_������ZS�#~��Gz���I�+���gǛ�tW�i3GǶe@M♡H�aD�(cڱ�M3ޒ��|��"�@S�jt�~�k�6��P
����I�����oZ�A�A�-��?e�1��$B��h]���/��31e�b8��R�Y���PK�O(�ʚC����������uI/{�H�f՚蔑g��-��ǿ��1�@�=j�b){�mxP���$oA�^���OXݖK򳥦�η;,o�������Ԣ��3��"Rt�g�������,H���pU�h�=�x66���Jg=��}�6#x,��8fl}	�Gy�����f���:�N�$�I��/|��Nn`j�62��ܨ�(q[���UL���3�]�V[̵���h���E���^����o�1���d1/�p�?9����b�*<�,�g$�P<cs3��Fg$�c���I���Vk�f|e8�F���?�C.ĵˆU6��O&�OZd�u��+!t��e<���^x��χ�/#oA r��6S���|��f�S`�-���q�-�! tq�@X�p���CB����$c���z�&Zh(��ǘ�Y�
х�9f[N�����w�j�8qy�6��G���>W+�Fs�<It��ܳ'E]h�KMy�[�ML��͖ �(�1��yhй	6��fD��$�S�L���j[��� ����[U)�&c"a���*���J��A,�+�U��u�S�D
7P�g�H����D<X�(5��	���ꫛũy����eDD���ꇹ!s�gws��ޮD����>��+��$�c�����6ȝle��t���A?ܛ�\���!����r��π5��f�?�Gwݝ�r(�z�U�-��`�e�����<���m���«b��x�m(�����'f�qr�C�!�!��K�<mj��L�[�deá��}�EQ�ȃ�=�_3����� �)(�5��O�e�4�h��A%���q
����Z����%����'Dn��/��Lt�M �R�-��T�8�N�ƞ+�ݮ$I�V����X{���КoL�H���~��p�av�w	`�m�*�܏Paqթ��"G8�'Ț�Z�|%��M@�Qy��ye�態Me�� f����[���$j4����^*��
"�E��z�y�5
�-�B��cE��s3{sq����5�#S��RO����~�`
��K�<�*�x�Yap\��f��ˣcL��2�/X�į�O�<��8�cBA�N�oJS=�A
���5~�_���se���ikK�Z��>k��JQCh��7�ǁ���鉅�e�Ju��x��F#�#�ҿ�Y��������� Wp�N��<�K�,d_�'pr)�P�ZŜ{DڼU�&���^`����K7?LUA�D�α��O��Jֲ����KH𙇜��tƘXkEf���3q�L�T��+��
�m&�`/��U���{�23H��]x�+����:���l�C���T����"���j߻~�@鰻~{�1�*�9L�p,k�~�} o"؂0c�.б��ëޞ4���HU�S}%���8k>�4:���x.�,���l@ui����fs�_�>�h�q��?��4OV��X�Q��M�Y6�p�)b�0�?�bFut��I��I��KwP=��b��S� 0��$��8&��<���Y�����G�!���`�QP�MUy�\8���@��ڿ\��t��#V�[�˱��&�u��5bnU)�1�p�L�c!����wƭ�{=��Av6���uȃ8��z�jP-�Y�|���y�x�	���M�[RĨ�o�	_,\��DX��|���ۑCIM�x���z��D� &h^�{L7�#���Q��U�� N��i�� P�^Io�f�a��N� ��R�7����U����:�`a����B�V����y�gm������ո:��c����ȃ!��`˥��ޱ?�3>�i3w+>�ǟ���%��� T_�+:�հOM*����5̥�!�6�Cl�&D�1��e��P,�'n�/ ��W�Y�V���~h]� ������s��h��9��4,��Sm��~E���bM��E���&⊎��$T�0M�P�0��j����h����@F |S`��nW#�3�'2�� ف���~&D4������۰r_�f��8�Y|.����X*�.fN�;��;0XŲ
sy
��a(�H���P��t@��P��
��_0��&0M�z��ƶ�mo+��Y��0��G�3�9�p���΀'&AJ�4�_�Yn~C��+���X���#��8�̰b;�����9*�VW��PQ�$ݹ��q�k�C�$5g���
�&�H,Ǧ��>�LE��1
!��ƍ��15�����z�g;���%�+ K�D1>�p���C�5�r�r��hu5�.�	�פ���-���j-1�x���ᢌ�5�RN�����0��- ¡���gƭ�Ŭ^W�K<��\.$\em|��9M��>)V�e�RK4Q�2�`�3^6���//Խ>$q׼�B�������r<�d`�L!x�W�|L��qG$vH�u���D��G�ۘ��
}g~
ѧ���o�:�����E-�V`�C&��`�Q߳Z�@�h�fY��w�we
�w4�Bd@�]\��tz�Ć,c�O��-I�b[��9����SӃ�ڃ�2�0����8x�]`Jȋ�t�$j�,m�-g��у���\F��2riM��uc�}�FS���w
�.�t;�Z��o�C�ӵ���0'Iɱ�U� �OZ�a|:�mִ�ï嘮��/�����|�KjN������'�v�!$�U�J�9�Ir=�v�*Z�d�
S*#3|Z���ĻB*��3�r���l��<�g�'�
U$�θ������'�j���~�!������R������LwD���0E�em��h������b��?���FJ��nЏO3�6�'B����@�j*��)�wJ+�ԡ���&-}���6UC����1eK��^�e$1�w�-Ci�~�p �y_�7C ���%�`�޴���2���u���G;8�s�h�xs�7/%�Z �.�?�f��ؾp4yt��YRFj��귽�Z�Ӎ��!f���NN�A��� =aXX������j�v$���hj����M`���
�qs�9"np�Ll"�Y�W%�It6�x��'b-*�.��ţ��ޮ�5)��.�.5Q*�J�q)kI��[>��ho`H-ꥵ5_j��F����7}2��Y:�n�ssp�u�%9v�G���e<O�k
�1�u�K�EG�`M�3������N0�ɢB���q_� �� ��s<[�Xc��|�Ip�Cf86�K��Bg�^��\bRN �2�g\����R2�wޣ�i(�K��,T��"U�`.�o�������&���6Xx�Ny&�b���A��8c.�S��73һD!(j�LЅ��97���a��[~��8.M�8̫���2�F�X棶�	(
J�$�]��YJi�-ŀЖ�فn�G���?:�PO�N~5ݢ3�;�ޚ��eX���T�cB�W�ejn��N��o7�)��$˴��'�Z�L��w�/�U�A�e�w��`���mGn�nL�=�1W���@.1 ��b�Kz14��/����<�<:7B���RN>�4 NIC�߲�|d�0J�c�4���'/b��\|ȡ��$l�3�$;Z�!g�K�b?�p�_�,5����)6�=���	\J���ޚBp��ƑV�#q 5@v
9_�|XU��Ky��	ɣ�,�K��Go��$��`i��7�^}�\*\��V��B�⅐����u�Ix��Y$�$~!�U�	�r����3	�l�_�"�F@�3��:�I��/��(Bfw#Α�q~�?Z����-����S�'�ʵ��8���)�v#��� )_��T����W�0�J:=-�9�8�ب���G�Ԥu�y�D3M�E���Ձ�t���_�Uyދ���`|��9�
��٤kՔ��b����w<�%-�@,�˯񀱞�b,9[e��|�-d�>�'Дf�I4ެ^�>��d�U��q'~H�^<Z4(��:��=��D	�]ȿ�#]?>�T8��	�$�8*�'���x��p���on9�z �)�B�'ki3����a���rl��6�2��N7rg94s��q�I/�/]����^��~�w�CT�Y�,�C�"S6F�HQ������W[�����(�Qe^Q8���*��#ȭ�8�1��Q��{��S�l��VM��(3C���F��>LI>��~\���aK�uLx5�GR�� ���C�FH9�]3a�G�/��xIy���1C��l)�v��c�3��Y0���fݙș�`�v�q��8@�	�L�0���t�(*Y?�g��p>�iO�����|i>|�=�A�nׁж�y�9��V#A*�QE�b{�놳�3.���&�ȱ<������>ŕTG󧇥'N)�M��þ{l¥�7Ȱg
��F$+@Q4V����q� 1қ��WV��j�I&n0�"ӱ/{|�;[-GAk��h#�Z|���`��o�
2n�n��Y�8i��GǦF�����E�؈�蝖G#5�EǩC-
��}�~zyC�;L��P����N����չ[S3jݦ����mR�?D�L�a�]ǒ��l3�}�5ȨGIJ���3N���P���M����c��0�%x�����"��U`<�{j�?T���g��o������c�}X����#ÜLû�MoBF�I�/p�V+z.���	0�u���]�^n��g�R
���aQi��$�.�mh�9�Gn��6�X��kX{E��N����֡؍���3���&*�xh㥈�y�G�6�� `e�>�V��[Q��5!��<b�%�U�\�Fy�$�\�l��ad����"�Q�W�ᆷ �9x(�E�B�­��?$�)}�*���t�tv�AyW����Q�yb;CtfZ�}5Z2!�c�y6�	U��?���e� b6�1���qntz$#�Fw�BN7�=�{�G�N�R�|� ��Sޕ�7o���9{*��Y��D����yuV+qjR!yh�%%ۄ�L�&�\���ˌ��j���yxK"F՚�f�*��Ӭ�d�Wkˁ|Ĩ.�˅ݡTW��߫�j��#����͜�-y�"q֩�Ѽl7`��o���ge�>jx�����N�m�7Y�{�G,�f��%�����W����z��Y�W�lPt�}�T���,�L\���w��e}Q���,E�;�a�=Z�"�Ca0�$��Ub�xcKY��Ҋ�E�8َ=;[ ��lڞJlړ��$��7p�k;;�&U��EK��ueju���$%Lb�%��_,s�o�N*���Պ*�����0��e}FZfR�F>�+�����|w�ΫHZ"-�Oe=.R�q��#��*�I�/�֊��s��2!j�O
i)С=�>o�&j��q�IxД<4�6����O>���:ۦ"�C��$�Zu ]*�!>�!���٠"$��W�>V���z��g�{���|��қ�� �K�q�8� �y�����y�l��A۵�.U��0��a[T���`S6�̎3���'�xݫ��!  �֠�ej���'�7��s&�y��m��R��h/5���gM��"���&W��K�v(wI��	#v�a=(�?�(�՟�����-����XB���b�L���@����)Bl������
�V��틀�Mۂw���?���¨z�-c���ȧ�nv�-޻�l�/�og�f���G�'oO+(���mI�n����|�c����]�Sve�#�&gr���𼌦���g����o��b=�4���y�|=RW�� �vAn�cQ7�2�E�3/b/�g�������W�� �1x��U;5�$�E�E�� `�]�;]A��o9�8I\4�)n\bmBBy�`���UI�p���yǺbA�6���bp�1��s_��Vm�{�a�/�&�
�AEX�s�h��'�8���d�5�(�$�i�$�̶��;ԟ��T_����|v�:]{�kf�\�w!ڰ�'P�fr��u9!�qX�eI}���J�0�a��Y�t�B�=d���|��a�b���g�.灅���YE���Ad��亂���f  � x�ـŐ�y�[��A%W��i���%S�9�ؑ�f}�_��Ï�r�6m*}=��7���&�	)m���>eg+�W�k�0�`�����TF|hS.y���d�A��/��!
���K+!Y`�_�V(x��h/۾�X�j~�v7��ˠ�C�Nd�?�>c��	�}W�����X��K�O���S�A`�1�Ɗ =&�-!�3E�kO(v�K��@���r�f<�~SaEN��T�O��Z��v��󟙮&��&��I��:"�c�a��=DȪJ�]��PC���[�LfX�z�{I{r��C]S
�F�{�<U7�6�>\�'���f}Ȗp����oȧ�A���/��B*�iH��"�8LUr?��DR y�y}�Z�z���l�pm.�
g��DpGc�I�Np�����0����"��r�
^�c`���Y_(e�`|�&=t=���v�ٚ����'q}$)�����s�\��D����N�	���#և���˱��+��~<V�=���lؑI��`�c�,e��L�F�B��ו�؎ �J�/�E����?�N�U�M��MU����d��?�=���nGB�mL��c�f����˂9I��O�'m�lڃez����_��1�\��X����b���r�<
���PT���� i���}X�S����Y�,+��7����)�:�\�5� V��N�g��?p��+B�3I�wn�7���:��N�e��{_'��*��zo+��ho��^����
����׫�1g�ii��ܐP8KlqZAZ�VG[��N��B:?.U6�B��'�U!�Nh3F~�
n"j�g�����gOU<�.������4���g���Uq�g뒂�W�F�!�)��'C�qO��6�t������p9�;ۊT�c�|e%���\�ӌo ՜�Q�ď����:Y$����-�T�`�n�!�6!ɒ�F��C/�|��P<�˫��8�;~�'�����א�˿�]	H�TL0���an8�є� N��u���H>h�b�Z��ټ?̏��;"L8Ie�u�6��u����3�Y�P�_�!�� ��
�a����"R%��TAL9�m�V;���B0^��)��Bu6�>~R�!H�T|�o�M�jr�����fhG�ΐT�z�2�%ѭ��>�b�i��m��J&������z�Ơe���Y�n\8@Tg#����s}T�v�g�R	�[��z2а|G�V{v�Tc���#���@Rav�~/V�0Ƽ��������N:>7rdW���C�	�B�gJ?T���..ك<|2M7�:���ߪ��g���Be�܏���F��e{rm�� 6qmO�3_����[r0���K��Ws�#���?)�^PNc.���.���d&R�� �;e�]_:=:���īƳL�B�V�rn!���)�ۥ1��i�.��<[F�a�R���C37<�,�r�jT�6l8%�C���G��ײ��� 1�؀��B��2P9�ѳگYh|�˶��4�1x-d����7L���x�0�B���Kk��K�l����+�4)��J<�r�[c�}"f��(�:Q/�
+�,�;ŧd�0�'zG�ݴ� �ǎ����R|���.�/h���LGX�vkz�Y��0�`I^N�k�u�>:=�3�}(�h���A��M!%������J�WI�hrZ�rMD��l}�V����
��K[ڄ:W�y��䴏�]��R��|p0�x�5��,�u.�ԁ��
A.�o-(�\�@K�Q��w�k�WJ�fk�s/�O��R����z�󳙏�6�M gJ�m*R�����V�ܔ�����D�~3��4ΛH9%p�^�<T���웎#��hb�s\��t�Z`^G�W	�����t�E���ݲ�G�p?�f�ń`SvC%ީA� B�~T&f,�|ź��W>9�ҤŃ�T�ɴ+ ��w���V��X�9�#���/����H���rCv��®���������is�%-�"�u]zxa|�K�æ�|Wʌa>�d#�S��O6���'!�u���9 �-�Ҫ��Q�9�rl��*~�#��3Y�oՃV���1��s��Z�5���c$��������fc���2��9Gu�[{`!�NX&R�ͦ��&��R2��d>^)�:���Q�W�;2���QR�O^���,�^ť"[9H��u~x������}��5Y�$N�������G�Hn�cH��W���gx���@�**�=�d�m�`�Vs�������3�h�o�|+�̗�T}��y������U��}e�w�/��O})�set��
9��%��6��"�y���Z��vO����AO���8�P�3?f������/lzƐ�/���X��i�p%�#W��1��M=o�	:���T(�
dB-�ޟ��;zw�2�&t�N��<ӧ@u^�2xBH�Yk��v��X�s[g�t�!���G0� �^�Xw����UN� �5�F�Ηw�Z-��^�^t�T`�I��rf��Zc��&^��1��c���8�U{?�%g���~|�?�!���l�:Om^��ɴ���ZdTt���z������&�U&�uҬ�㹊�{d��G�w<G�Iz���><�����k���ӅN���E\ͳ|c�e��2������6�YfLm�"a���8}u�����d��W���I�W�>�}�'sÑ��Vq��D�z�m��׍�*�*��}�ri�D ��W�*^�����P.Yt�y�ݍOK�e���"�AĖ
n�G���x����/��G��.��TT���wXR�җ2'�s<��eVw��Ş�%�(B���"K����LxGZ\jRt!Ld� �xź-K�I(��-�����_�Lω�,g0��u!5�x�qC����$��<8R���Ԉ,�'B��"Uܽ�R�K���՜H��?#(���8���h�y�Y�4Щ�7M��jfM������+U���9�����8lf9V�Q��3Z�v�r|��x��I��/-�SkCnz`�������LF��ׅ�O�3�(�q�cq����1�Ȭ�\�3[�"� �[.�z����M�5}�S��'JxIUx��8ɉx����i�Z9�z�jR��\���#�nƓ���U$��tbH3s��^!>Z��=���ru3��0��J8�$��:0MOS��'L'�H�%����b��������\�+s5ɡ���C=����Ρ�-.Z�	���U�՞�ok�*VƷԥ4`l�'S־N%,�8����G.xF&����7⥗�&l4��_�ſ�"n��g�oZ�\��=$3���@L*�X��ӡ`��\U��	=��\*�����:��@����f��sD�Ә ��=dk>��YqMiz�G��7w���Q��L���h����/���}�/,�>F��g�U(܅n�����bSʡ�\��utv{����^� c���P�����_�	�|�!�!g�#�f�ߦE��T.d���?�41'h����q
���=���`��h����jl�GnN�����+�lB��Q
S�*N���Y�M�iK���� ֮����'���c�X�j�K�Xh_d�5�u�>gJ�
�t�`�t�����pPX��lc��Y�g�%��9A��0��W=��\؏^'���yA���1�����Zb��8@d������J����������M�1�+k���#���os *�aR����qXX��} ��w�#���9x����U#��(���f:ve�e��#L�����}#���x�9�I%�b�!Q/�_׈R��d�*O^��/��֩p����_l�\͝-�`�6U]��_M�ϙe���c.B-�`�K1�ZXg�Dm�Җ'����������y�F�`�F� P3��)�k��ͦ�k�Ǖf������
�~(s��@wi�i �Z��]$A�B��������}��������2�@�õ���ٝ�O�S��]!-j��{�W��-l����]�Q׎��<�Ȧw>�2=J�ɤ�v����0ˮ�g�"�*�_7?E�0FՆ�J��ϭ�qal�̸"��>�8Ȑ8>��%Ƽ�!�A,��7�0�.z�s�*=ӮL�]]7��ٍHPaCn�p�<4�qw��폹�U�s���_Bo]V�l8���,-��U(X��:.1��TA�i��X��I[��i<����I1nCt~c����
E��9E8���G}-���kߑ^VD"���"h|��3_4�9._@iJ�Eoӏ"�����б��,$9���VO�XW���/B���Xg��$�V�09��q1AtR��������#�s�s����^�q�2�''�3��˭|�ϯcq�gDb��8�=<�A<�tB�.Of�����I3��,l��sw�|�@��ż�rH{����&���k���k�
&�W� U���H���J��g�n��ԱX�Wrl�"ꐍ�1�_��^ÊK�~�_��qn��_�]�+��u�������6�UGV�wN0�U�r��  Uz�%I��R��6�X�0c�n����X���78ui���Fy�t��~^��g�)?n#Ʃ��oI�m���s[����& �)3Ooۻ����Ax��W�gczQ �>��66��д,si���m��?}���N�h�0�R�o2<6�>.���_�48b��wR�Y�9��t�IQ�t^ˡ��/��=�C�qX�A��R'�g1�����ԍB��6Z ���H�d�������V�r���v9�u�Djw��Q���n���QqV	>S�'��^��k8�9j����S�(`���R 'J�2�L�P쾴B��?�@m�C�#;��(7�D�a�v�N�@�>l�D��\����� gZe�7Vw�>E�	UZ d�Kٴ�@���f���}��Z�$�;�oh�����6Ѕ�$�j+R��:R'#�e;�f����������CZ�@�t �e��@��4��{�a/�P3]���9SW$�I�8fTU�t}	4�"�%��ߪ����XMJ���4G��N��W�Gq*>�o��JJ�#O�c�($3y��D�>Vƾ$���QP�'�m*ES`�}"�}r���nt��UV�F̸�k����PtY7�}0#,h;�P�����:�^��ǂ$����Nh"�������/�Z�#�Q��C�S���2��!�i��@}�z�4`y��ٖ�H�r�}7����i%6�T�Duz/��c�:j�?I����Y3qmCM�z���tv��h{ ����39d���*C��Ua;h&�����h�-UP��pz���E�g9�u�|P�ϝg�]���.
��Wؙ&��L������DlC_��+����}�P���l����B�;Xk�/�۝�p6~�T&�H��!*{>e!����cG���zI��Z���9Y&<ٯ�^�2�bI�c�9�
d����њ�Y6�@��s�R}n��4t�O����j��)�M�72�q�f��j�~���4S��·�ZZ�b���K��ڎS8�=���@:FH0f��	u��HM����U��P.��q�"�g��U���QIg}�Z=J��H��1��ǳ�����ُPj���7��g�����mݚ;s}�'1�3d������\�螽�D��)�Y��q?�ڍ�+��ݾ���BuB�3c�Hae�"�E_��3��k�8��a_��d�c{�5r�\��C9��:D��/<\���!���b�4WS�eB����զN����z���R�������I�F#�p���B	�F`�X*��\��k(Pg������M�T���(/&0W�	{lq��@�y����<�Z�[�+6i�V���j��#1��n��j�e��d�W�
y��״�N�"q�y�ӎf���"/��mDo@,�i~���к��~��#����bk�(Q"o0/�[%�%�9�j��oaP�-">Χ2���H�y�8�U%���D�&���$x�(�_����i�U�ʴ�UDJS�W�D�n4�5E�3� fD<3Pw>�s��|:^_F�%R�hXrv@�)�O�\�Z���!()b�D�:��[��6f�o�T�f�$����>;Ji��@|[�_�kFC��\�T5�5�v}e$�kw|���J<�;Q�BS���a���QN��taQ�C�FvnY��E7LkS��o���(i�w�Tz�Ou��naT�15�^�3؍�(�)
A|���τ�*gSd�[.�5kaې��eV*ro�������)(�q2���R9�ʭ1��:�$6�}L������C�(I�\�����ov�m�Si�����T-4�?�]t���Nz�"&WY+��&�Q�&c��Ѱ!�����I��,Z�]���FSjJ��BEZc64�ul���j�,=A��Ux59���&H�qU�u)NLut(U̕M�h/�p�����q����v��)�^�w{(=�	(ބh�H(�`s8�QzJ����ám/Ǵ]�:����mY(YR���!�ծhlCB(�q�L:mmVnT�=�������D������l�1l�H2������^ R�JoL��
���蹉��y6�;�����A:�zP��������H�� Qӿ���,�%��x�]j��^ѿ�B$��fT�P�wiEJ4�-��(��Ֆ"�r��P�/,�J']�$��,Z��� ����ېkr�=�("�#���݂EnƸ�[��1���p@�>����Qѣ�<����]����D�mC8S,�V�?�ݧ��f[[�L��_�![���m�lI�z��-�KQ�"5���kʣ��]y�d�Y�x��? �V�P������wVEI�M����Z���fm�����ç����m�0�V�{��=��A���MN�]�#8|����x�I{q�ZAa�u�*Dj�ù�	O����'�-_�@��
��<�(���ǂ�g�!���[��즵��������'����2�l�=<���yl�mި�諎B��w����Qޮy���������N����H9����� r�{�d�.���$��Td`��g�-A˙�$ǌ���ځ�^#������ I�
�?�ؗ��O��
н�~U�_�)�3�����u��	�A��А-��]��Ġ����O�U�GF��@�ה�m��?��(n>�錪�ktq�𱔠�cuh��'��{�pƚ��<�8��~�����f�N�&ÒXe�R�Kqe�:K.�Ǐ�*�O%N(���y��L~��֛�Ҕ�Kk��n��`㘒��2r5�{=\�D��9 �'w��SF��]<<зq��9����0�֢[�p������<X{�rcr���_���i���"�Y:`I��f3|��\>x��9��O��-�����xUM�_}n��=�����m��T
M�v��%���S@(vz��np�������9�
{����]��?^�@W�7���������@Ɇ`�]�Z�AtS�nG�H:^D:VW�A���ق���Ȋ|��Ѭ-�	>9P �Э'�+l��W�y���n���>����L�*k;�mOUl!��xe܅��e_Y� �Ւ��3A2ܐҙ�"Ӣ)��{�i���N�����v�#*n����}���at��碽T���e"@Qj�Or�O��8���0,*aM����o��*!(������ q�����P�Sp߲5����� J������5��0�ǈ=洴�]�vj|.������<��sO�iH;2{ST�B<�����FM��7�H�]��}i�ݾ{�O�<�D��i��LZ��p�e8��pz�i�Y��&w�a�����6{f���������Z���Ƙ��g�\�!�WC��ӏJ�[�"��Ҷ�k���Sh_P��7v�8k��\�uG�C�Z�	?A��4�}eh�ьiiO����>j��6�}h�51U��>��l5x�-�g����k$J�p~W��
Z��-srn����� �8���#gWn�-	=z�î0��j�����1�s@�ޟ֘����(�<v�`�&F흋u��=PU�,���q�w5R��%�K��-�H��*ީ�I��Z�v��U�"*���k���x[2�l>�x�H��Gm7ܮ��5	.��u��b#��/�&Y\�(A���zC�D�q�>e4e�� j�׵Es��[�sql�(}��Q�[*��Gp��H7�	�@�V굮�I��@;�]0�\)� �7��joy�OK"�Z�Y��@ ��T���_��DP+�pQ���s����fc�XR�yoD�_��]�U�͘�3o�FŮ�ϥ�����©Y��H��)2��_�P��5��J"O�c��f�����������a���2��n�	�N��/��M�RB�f}-~TPܖ�Dai^cn#�mo�����`<�_!e�zC�V��I>i"6���Eo�}�T�J����8N�Ur��1�D��������R���ݮ-��sq�hpGEi��1(�:��sw|{g��mC($�j��2ݡ@ �~�wWٜz����d!m�M�Vvo�h|"��#S��$	���}���'��0tL��l��Wᗪ��2��L{ￎ}><�)�����U|��B=��JP���ۣ"DOKh 3!"���H]\gBI�SP])��Ė��7���$��AaFR�ڃ�7�,J��9xmN9&e<|b����Éc���Dc|�.ט�T�<v��G�z^3ϖ���5������"�ڷҁ�L�5��H�Ӯԁ��9oW���c:f��J�0�ƉfN�v�\�N����}�p%>��q���.^��9�l���s:E�x�%v#��bՁ��L��`<ǍƘ�K�^ƓJ2�L��)3�:�<��s�%b|u^�OZ}��p(��E� c�ܜ�KMCeFGۍ�*��>���f�/[��m�R�K��4�-��f�bsדP�ě?H]q�{��ڤ^i�|5�C���S��f��b=9�%��Aa��'J�Io�@_``/N�7F�,�\�S�:�ܲ>neL�z����=M#:�q4� ��9�KgEY���n��\N�+"ڣ��#C!,���Vo��s|kժ�U� ��K��e�W(ne�������G��O�������']<��U�_	���9���z��������Tɬ�Ċ���k"J�3���A:n����M|�o���*O��I��?/�Fp��b ��S
��ˈ�����ӹz����-}�yx�d�G�� )���� +�� ����]��Î6�-)�74��9dd1G���9�����XS�7��.����4ld����o5]�@`1?6Un@k����TW�"�|������j��Sڙm[�
�qo_(?�%h6 #�%�Ɍ�S�I|4���$PnrQ��	�����x_��WRr�>��,����s{��/�	�q���T�¼��������C�N4�C#	~��`ܮ�b1����c�6��__�gl5�,�]mZ��"���d�P���ą
�5��>�����;UkLF�����i�K�T����&�bCw/Չ��V6� W<�Y�KI���j<�=�f?�ɠ����`oVP[
���T��X��+μ��o!�[6F�bA2f���g�2H3dY���x�M�ɘ�s�ق�9��W�fV���"�7��6Lݿ "�3�bUO�ٛ��'��˾ݾ5�Tq�sS�3��-N�8��]�@���E�ˮe�A���V����pr�B�S~G?N3�Y�nn��t��U>�̂;��x(��mw	|��/�3Mud��i�z��
�e�JW��ͯsS�m���V"Z�����D�t:��7�G�G�ʤ�;2c�T_b�s�	���M��؊e�%��O����5����t�c��h�\?/b8�H�eچW����Hxڔ=6�5fL-ʩ6�
a{��k��(�zM���F6=��\��9>")����ԻsP1Zj@sm��Y?��{a��KU���^�dH)Z���"���1ʮR�&�_�,��T�ak��+��,�$}zCU�S�Eo�u`}�,���-_L~g GP�{*n���~��W�V�5�3X��~���j��?���������ȩ2��!���)�p4�w�7���I澌�,[�i���]�k?��WāU�y�n�"S�R�D��f$�a�Ғ��Y�>@���(���v�n>*p��H/j�| /����*r�ADI$�+���t�Յ�7K�ݟkA�9��z�լ�4����=!���?�t�L�ig`Pӣ��6��*����|�q���a���|/s�t��'z8�V��%�uæ�
mE��C|I�D���~��gh�@���(һ���11	.��6?��j54�dL���Ð�M��7��h:��F�AS!��پ�cd��)���Y��^�aջFe٭>�B�	{]��J���]?K{�juK�>�Fl���W4|�0�M�wI�aƆ�vN4H`/@�i�8�%A����S���ں��=��v� �߈�49�?%�C�Y��!G��9� ��E*�R�N��� {�t�N��E��2�=�{����<��Sj8"(0�2�`��?�G	(/�˚��[�g���~M�wi�l���Y�-�7���I�OP$��x�->>Ϋ�re{6E����>r�p���?`�	I񘙚��C�%R%!��Z��ǧz�N�bD���Z��ݙ��j!�1s��ysJP�v={m*� ����_����ib�>�>���xs�b��)P���)�"�z�V�|D
A� ��e�_������
�q%�H�E��'����`�����.e:ȩ4�B� ��@��-/���	�,0�n�Eu�z���͘�ʙL���R]6���j�q�Uc����|�AjŀWb^W[�-V���8��R��_f����+��x�~��R����C�VR����X����[c��U{P�>�A�scS����O�FO�ʗ��� �o-��a�q��C���;��>=F���"1��i�V���Ʃg�\d���Յ�|�v�-�|eu�sط�d���RU�����Fg��.����'U����2&B&�Ŝ��ES���&��86�JҧŕxvɁ��
�o?li�\�>�A�1t�О�v��ךal��Ձe�x�Uu��K���
5�ʦX��������ް�Rx�'�!�S^J� fM*m��L�:�i�*:�\ ��� �����q�hÎ4�6$|�gl(�{�rה�T���_�Sln@=�{y�9	@PA�l|4gbjnt���5��v��t��d�3��A ��5DL�d��ƁP��
����<�o�8�qBɉ��"7��߶�)��]7:�a��2Q��3:�� ���xQ��'��ЯN�H��xc�f0��C]R����b9'v���d`��*����z1܎
�����(zRޏ�Wkn)5%)�!�1ͻ\a�7TPkm�n͡R
7�wIC� ��AF���Vy��ζ1iu�yV_i����&�B��yDadW5�)�VD���E�ZжI���A�"�"�����c��@mv[���4Ͷ�D�@�'Zx��#��V�Y>�xc,��Y��B0R�i�E�՛$��{o�� U��Bߒo���^����`��^�kǴ�����#j5/��D%w$��.��L.R�+Gat3z�����&��Zb��T��Z^���.��o���C�"C�}�hє'��Ùf��%��	F�mb��ټvA��x���B���o1(7�;^�>?��f'^L�fJ���^����[	�ԗz�:�O��x8��ӂdRXZ�kż���QU$B�-�"C�Ve���j��Hm�>����)�|Fr�T�B֔���EXw�b�i!o����_���
�ި����b�䷴��sW�p�EK!���I�4��8�LǬ�KL[�/
[��N�1 0J
��E�ީG��J��g����o��!���2�� !��o*5��C�.��@ҁ,�a�_�M�+qo7$�j�����f��0��(魱��v2s���.K�J����jR��Ӕ&�,��Ę^� ��������؆[���?��\b�U%�a㎿U�2`�&�A���L��7��[�,_��/ͪJl��ҁ�N"A��*몬�9.!���'�X�F;mi�8L�*�_��
�<���xS��� �X��[R���c��U��"XD�;��0���u��a�%Zu
���K���5�r�r3�fl-IVW�;�{�$�k7k�w���	|J�N0�f��9���e<�3��ek�"���ao"��y~�qMȐJ���2�|
��T��e43��q�h�ɀ R�tu�v�:�4	gao���)=L��=í_ۆ1ˑ��5T��e.hƑ8�*��߁��[�3o|�^���J	���u���[�^0cv0һ�4�1r]w��<\m &/5�[H�<��HǶ-0XB$��C34�<�-Jɓ�h��/��H^�8�6�����7����}9P�	�.��m������=�#�W�M���{@��)�����2�t�u,�\�픏,�|�=�!ˆ�.P}�y���˚f:ۓ9�X�=�1�������\�=�?�� >����g��N��-��Ӛ���d�o�	��F����w�}�@��Ba��fk	[����V�,	�z���L�1!�hz{�M����<��y�ڱ�� (	i��Ϛ�~�Oۗ(��|��T��9�&i'p;�Ή�E���V=VYp+��x���%�O]���@D;�b�����%8%&G�ըW�'g ����i_�)]����F-��t*��� I٭h
�J���B�� �t����Zk3�NA�F��u�ed���n�E`�,=6�����a������t�Z��5ˎ�m��a��ڮ�jw��X�4e���np䴛 ���';��,q�K��q�謟�([HBЉ�7�c�����x�to*�>v�i�)�?vd�۹��ޅ<��7Pj�X�Sj-)���Yӓ���$��V,)u���m���1"��C�؟����r�eL|����	���?2z�6�F���+,�N���˂HR�QFA���� N���B8]�.rt&0��1��z����1��Șd%�l�_�[��4�fcV��]����qHhD ��U[��:�&(�P3�6�Х<x`N��������&��yTM�'�R���HןVhA)���D>�	�o�F䃡��ne\͙�>���:�{�AX�sj���8�m�o2YBB����ݟ�-L�3л��"׈�3Y$����<��������lg~��fJ^���{�QƘ�j���gx�V�j�f�[����?1]���F�+��8�t�������iaа�!��M�a^�[	�G�j��SCE�7允��^��=;�����K�}�
G:���~_�l؆{���I�w�$�_���t4H�m��eJB�t���b���a>E����J��`Kl����ky���w�>$$�ِ���������e��G �s���i���M�ٷo
@��V�f�J��,̕]��x�lFmL�����=!� �d)d-����j���Y�o�6Z]���./d���@,z�7 �XZ��т@�ZEr�q�f�����#=��ML�y�~�V>��7,��u26m�(1no
������2A�H��'�����$�i�%��6I9Y
X���ٻ�WU|䫣��G���d 咜����� �tַ$k{�)_�?���ӵ���	�;�ۙ ���0p.[��:�#��,Q`�IZ��O�{YD/����^)8@d�'�&OJ}�j��>����~er5��\?u�h�l1��}�DQ���њ�/"���1m?�A,���x)��m<����7k�iH9 ��c0����+g�<bA�4i�qJ��5�Oj+�5��avj}xi2�C��^X���6�)N% S�@�r���&0�Y6������wb�Cx
�o۶�[%��-��&^U�Ey�ʺ����I��<K(�r��?o8z5�i��P����_��c��ηлz`n��ܫ�Gʈ�`��sZ7�o��=E�����ٶ����:�Br�K�\�z�⁎A�*�-/�/-��������h=+�e���Ak�1uU��@�.;E��MB�q�מR�T���2��<dF��H��Fe��^A7<��K2h������+O.��*�F�3���+�
��0�����q%���4�aМ��ts�@Gn�ܹίO�v�a� �w���)�)�W'����XDe1�X.r�ņ�k�M��8��wf!u���m�-��9�N]���~<���ڒ��]\�ۃ�h���4��;.tϞX�j�ǚ>F�/sN
I�i���F��Ӧ{�̴�Z����]���P6j�&�c�͊�}X�d{���t'JD�}T5]+B��ˆ����q�`8���/%K�u�J�N�ٚ�r����V!UZ�i�Cܡ����8Y�m�Rԑ���u��y�s�\]�`H��K7�.��	g����>8�+}�L��"�6�,ox�������������_O\�ʘq:���I?���5���{9;�6(�x<E@��Z0�KX|�}�G�����F�ԛ�q-*�婰��&���i�3z�w����թ\�56tdC=!�!�!�HL�[%��y�D�}46�3�r��V��<NP���3�t�1���=���0�n]�����?X�M#���0�[iX�_��Q<���:��ʊlq=����i���,�� ��9r��Uף�u4?��	����:[�{��X������݀дZ",�6�W�c����6���3��W�Nȧ@]ڭnG["�s� Dv���yp�8k�@�����Lw�Xc+ X���<�=�X ��f�������`�a����=%?�G���n�⨍lE��~h����l���)�R��~ �le���Y��Xw¿s��u5h����b�-f�,�����{�H�i�������)y���dk[�=QU��|o�s?��9��1��WV�Pc�麳��VS�7�R��40��Χ�|R�rz��t��:���	t+#I�3�t���om��>9=F��0��@�H=�����	*g�a�z9`!e/�>��a�X��Y�Bn�]��V�#1��l�W�m�Rq�I��O��'�0г8���,Uю��6��Ev-��/F��ɼW>_F��yȏ����
����{�T��	*�r�0Paxf��9�&��%���r,j.;�R��x9�X��d��2590�UF�{��g�����:C�^I�wKG!��/O�6��$�OqB�Ս����;�V�KU�뀺U�(P,�s�����a�ǟ=og�����cT���#���YH�6;���K�.��+\Ҫ�ͩX��>����2��a�~����`q]�̞����7?���rX�/#�D/⬒��]0�$S&,��,2l;���k���.¤:�o^�)az��.1e
�r�E��A�Q�S�5&� ]�<�h[��i��$�@�����#�պ�g�=|m�}�����	�Ĝiu��l{m0�H#́t��PP��u��[8H ����C������*�/Ś3�/�`�6�l>���2��o��L�W��*�Ӧ��w�6D��[�C�m��ߖ�	�I�D���Z����3d	�IH�1;c���8}�4��g�?�pnnZ95`pi�d�UT _r��XM�)��6z��֑%�������|hK�z�7�~?S���F��������1Ӣ	u!��B�2����ދ��,U���}B��H�(���(���ls�;�C�reU�� ]��?��sv0f�-�4�w·a��ߗ{L��N-��WÈ� ���An���M�bRZ}E�Ԫ�P�u��:�:+���&f��D�W�He��{�nfSAux��!4��V7�^�G����Q��q:�W&OSa�s��i_����~�L	��Kh[1�B����AR��E�(�,�C��CV��25fk���	4{�q���/���c��=8	>z�f;p��d���˯VM�8}9��M'A�Se�0�輬�:mBf�@J�wT�+���Ofh���o����������M�[�:v�R��9��1b��������������֛�*�O��Hd�`g�a�m [ɷ����������B7}��saD��B������&.���wԑa�/��*���Kj�VL˷�)�-G��)x��b!HcU
�}��A9���4#f;<�@ы��(!@|A�qJ_���5�r�>k�Ԓ>%q �gK���`��nJ~O�	Rz�;@��Xz'}I�ج�;)O'��'f����aZ5���e�S����&f���7���@v���P�x�پ�O�_��v$p4{���}j�d�(�k�cE><z�f��z�J��)�qq'����&�$�޹�8�~hO�>�J8�St'Sf��N?C)�Z{X'?d#�����3���JS6��0�/���6�kq쪤�E�r`!4�w��'�=����6��Be�����S�<Yk�4-Aq��,s���YH���wv�,6������4���v���f�.�J�^q*|����#�ב�+U-��tD�X,��.hq?z�)���:s��#�Q+���V�о�W/5r	��iޖ��'��m�"a�.��s�����g�ӕJi KQ�W� �{��V*q)�WN!�c�����`W��M��*�^FT;rt8���\���bAz�H���s��i����aݑcPL!A��릲	�Nwf��0�X��)=��.Pk�����Dĺ~&ɛ����Ns�hр�vz1L�#G���F6��H �d���c����/J�ۄ�ޙP)ɛ�ቷ�G�z�s,aDg]K�σ_3�;\�6��fi��Q��1����'��2����%a�MG�S�H����L�pY�|����RHcɫ����.��gAR���{Z.��/O�i��m���v5]j���\?����Q*�6cipr������ͣjS���	}���γ���C����k$$�~�M�x���,J�����.�cX����3�0���"t�ޞ�lx�G>�'ѢsArS��]ȡ5KSB]��<y�˸�K�3S9�q�P�j�Õ��3�����+n3�tl�Ru��Z��d�B���t����9���'��)5r�h���-"1Z,�'l��k#��t13�U���W7��
0�Vד#�O2���(��Ļ:!#��_
�.p�I���I��⒨�Y�߹��OHQ��O�%�&�.p���u-��ј�Y���Ȱ<�~���$-ۛK��'iK�|h�O���7;G�ْުfϙ/G��#��#clr)FoU�&$"���*G�"�3w��%�F'�{S�^QM��`s�۩,�����+H���%�B�:��/�F뤅�Xs�)�� D1,��#o�W\R������'��X�[x(�ȥ@Ts�I�ɭ�kAM��_2�2����j.��;�Gc(�	x��H:��4��vL��'�J���BFH��~����$_���m�BP��Ʌ7^M���u��!Z�J����E 3�-L��-�*?r�E�'z�|��#�^�K��I��|����V0�V�U	%(f����;O��C�!z7ָ������t���i*!̌ �OVXd/^�Z��?�����������1���R�d2�K�iH�Y�HPht���P�&u������3�m9��BK�d:�� 	��Gv�E^dU�l�����63��u&Uo�$|�d@��n��^޷�)����4h��������	(�?v՝,_��y �|vd��·��N�J�D��zgi�5�"��]}�ĈR���� ϰ�I����@����4�%[�|ܿz��(eaPW#Ha��MIW��QCb0=ae7v�f�g�?)d���Q(���Ni�`r��0⸨����I��aR,t��
�'bJ?e�L�{�}��������e�y��m�7��WAe��-�u�6�	
�m�x7n=lEW��<�eޝ8���dզ- ��ysn
FCU�(0��5j`a����=��:D����|�z]�m������E���A�v��3��~X�9@�v�{<`�̍�a�hDƍ�&�ڔ	��X5��nMH�C��<����#!�d���@�ye)����B�� �,��VGx�}�0*1u�ݤ%_��d��(��Q�~�i���@��4�ش��\G��u�w_44�:�iw�M�1�x��rt٬LNQ�eI�7O�$W蚗N���)L�09�7t̺�m ��i�.<�l�)����ۤ��Y�������X���gfl'L�[g)J/8ɵˬ�;m�K�
�a�G&$�R#,&�O�e�ƁhS �ø!D� ������D1���m�{�b�L7�PƴtWYKcm�B�!� l�t����l��x9�U#{.�;xi��	��7�ҏ��ծ�4�p����E�FŐ~� g�%w�h}Ɨ�Gs�>�q�h�٧�b�S޲'�+��r��u�P��]s�fd����|�s�'����u��v�ՒI�����?�|y��j���F��LR���u��}NϋHs������?<zo��d��2���k�i���a�˕�K��(��L��8�у%d�9��jC��ܰl0i���S}m1�5��'U0;�������w��IB��T�[l�'�-��)5���<�^��j�>�.�2�E�gP�5�'�����%����Q�(~
L�r��O�� 8�M��B=s���s��j�Y�0�_%�omzm�{�D �(���Μ:m��_QȄ#.Lʗ�N2*U3����=;ߣ���
�FIԔ�ȗ���YF��2FX�S�����T����7��
6�n\���&K��K�+���8t޼�Y������X���M��&��8��ު�~�1D�<��0 ��d6�z�͐w��=���I��z#�_�� ^��ܳ��K�kϲJ1��QoMb�(ߝ��s'U�Um��yfv(g�P�*m�D=���>�N�۠�5>�M�����IO:��-RCuG�~8�П�#�����fX�8���A��V�z�����*�iѶ�11��/����d8s�c��$�dM��7M�63��b�c�;P)�4<J%����2#�8(���Y�4�W FA�1 �I�&�&�U^��ĕ���,%���Գ^c����bt��ЩQ�6�ϛ���WE��>'ĒfFW�a:J �L�����×F=X�D��0B�u�n!��5	lBW`�� ,7,g`:	�c�EJ57V�pO�n�nq�;3�2���(:OJi�ԗX��֒!���Yp	�{N����EM�� ��7k;v�U ��.R�k����2���p��R"��X\��2��D���q�K�ʏ��|J�A:�}��'�x����*�;����k��?V�����v,��g�M�'O��Z�F�RFT'�m�������I��ihg�q�eŴW�5Q�'���h���t�˅;[�ߝYk�+?�V���N�g��n��7u΍���S����#�ܦ�A=�cM�`�K]���Z�ua��Y�p�0]G�F�r0���8��c�f�z_$N����'E�׀W�
]T�3eHO,Yi&@�(�3����~����.��U
g��_���b.<jDǇ?5�>6�~���_�* h��_܍6h�OB��`�PQq�[�@L�$5h��x�@P6�k ��d;&���no�a}��:�2W�k��X~Ri��f��`��G\cD�w���or��	CBF~e�4��"L��#@!�$�ǌj�j DL����҅Mf��ϗ��	�4�"���ʚݷ�8��j�Iq"��Ծ�!$�h۞�O E"D�;�kňN"%(�kk�G�� `s.$�0�!��)n��E�$f��{�47i�ا�X�m^UM$�F` ��4�闰�+�(�ɋ��O�!��RrG�6[�-Q���)���6��9&�����0�.TZDu�K���_c�#��)�{M�~�g�OL�q��)�� 	�9��vJq�_�a&�q��\�B^�:E�h~E�J���-��<=C�%6R�a'������a$J���Ut���Mu��6E�	��$H͑# �bzˆ�K|��jA����#(�KZ>��+�S�j�q��)֔�+?`-i�l��~���庺"���_�������QK�(�G���ଋ�ø���=!�Q3�F�����\�<�	d��b��m��>T��{��(F��У����S�0�r¤���]C"��,����p6K��MA��P�Ĉ�TK��]UT���=�+y�*�1�3f�L\�==Ά<%܏&����DT$�F�U��*dxb��q�IHQ���Q�U������ă����w������0�W��|�#Jiыj%�}U����k3M��X��zn)
8�<
��564e� 0Г=
y�%৅��-�EP8�	f~H�X����?Ȣ�KU=D��|���)�Yj=��R":ks�h�y�Rp�B��T�|�VѾ����tg����6"���ɜ����PZ՜
 �t�8�=�-�AHE�$��X7� "��L����AҴ65�*��n[IV7蕜֗��ϖx;�S���/s�L)�"���q�o�T�H���[�艾�������E�(d�8Y)��aL�Z 8Tj�P�c{|a����|XT�P��i啌g#U�ѷ�)�_h"��:;q�
[c���c���+r�ke/����'+����|I�:�'��UۗBU̠x%rX���ﵯO��H��<D��ʟCj=l�{_^�Z.) p\��� ��cܑ�]X/�[����}F%~����z�3�& �f!%%�޵��?yL�o�4\�����?&�k�4�8Ny":����w{]���٭���?5 {���mW���8�6>j�|�G)�I�ް׮�ߒ�>���H�Hw�=���Zy�~8��;K9ۯs���q�p��	��X�Ek���RL���ۆ��!l1ݽ6j8Y�[����_��W�y��3�98��"|���|�_
��D~Z
�L�Ɛ�8w0*� �*�t����g�n=o��uX��|<x���=�ct����F�D�s'�08T�у4��&T�S�pW�{6<���@�b<�GǕFh��|��[B?��F�蓚�� T���t�n���9�DҎE��ŶvJg�a��u�Q�E &򗃁�Gy\N�諕A��d��~�ܺ�i�j@:�2�GZ
�T�� $k=�C��&E�d�PVE	��!+�c���a\&���'$��G��Y������*(hÎ���ȧ
ܸ��mJ�Ψ�����<��5J�ߢ9ta�-�N��V�=A�خ��r�9�C=��a��jZ=��ú9Ul��;���*$�B/eH��׷˅̙� CP�>o1k{~3%J��p��tt���,V��@���C��B{7�ːP�Ǩa
�6�pT�:G�㉑_��z?"\�� ��V���G�E�W+�)A�)sϝ�o{x=z_4�^.@��b��B������c�}������h��f3�F{;6yƳ�{�M�p���؉�|S"@#���R�~���oK�|6ܙ~� l���k��O��"��Z�1����s>/��7���(�T��� ݘ
�_`�ׯ}V�@ȥ(a�=�'�Ej�����G;��؉>�tp��D���4�4w7�@�Nnn��%p�wyQvo� ����!O77e��j/���{=�WRb�u}M	��O.!� �܃f�Τ+S��J�F�X!�e(�R[F&�]8ج*1wR.b���lfQ�Dg �M�HQ������O��:�Ci>{�h������Ey��>�Xa���[V;���8�+�)�1�	3��H�k|C�����Ȁ�Ҁ:�r�v	�bS���\U^Ӑ��X��9n,�Q]w�����N�I n�y�[)��������!����i
-����Ĥ9ʸIe�R��=c� S�CMh07�o�f'-6g�]ͅ\pC,*���<�P<]e_K*��Ŋ%?�kH�E�je�q��z���!A&`���mrCn�іߡ"b���*��Un�_�ǈ�Fɧ���f�,������
��ٵ�n.��&_��*o
D[�L�E��3�h�S���י�^�����xZ��h2�*S�YP�D�*�ǄӇ6*����"�,��<+*�~�DP&jN;��hHQ���/�{��ŴW��`j��GޡJsշy�uZ*��;&��Զ���F�����ˈͧ���dQ��痣M�PTL<`~���ZNV��pr����K���Ow�5�]銌{����Bf�Fv��w��n�ř1�8��b�r:���뭨C�>��K��f݉TEW}�cFC+�niى�u'�bk��e�W�L�W��Mq�[�@B�����d%�L+!��b��B=h��_�Ӕfsݕ�sSI��{@�G�#�h�@2ը�R����\��K=����"@���{΂�,����-�vN�-ϐ�@�&���_߲��n�Fȇ��.X��"k��8f�C���~8�aiQ$ ��4w��J�U�S���xʾ�� q\���"�^�$1�<�����	݌�W#�.�7���yP�:0tְ'���Nذh�Wĭ��YG3)������&�[8�IO�O� ����F-1��Ķz.V��oL2
!�B�֫���'�S���UM���@F�����(��:����yb���������#�K� }�=�x�<���g-t<h����8���s�����:�ŴLr�����BOʮ�%|�ڽ�_[�!��RlA�l�ߜ��AҎШBċFr������;��B����J��M��Eb��iI<>�h"�a
��ݑm+ �v��@���a�<+�]^"C.�8�l6!����HQ;�$�s�˾�h�(�d�jP��GJJ��	$F���<��ɣ*>��qS�)���P����e{����9G섮F��=G���a�Q��Ut�t�ܭ^KO�}ը����WvR�y<�E�uQ8W���{�|'�?X:T����7a�%�Q���n���r;�Ǜ�H�� ��j��&斆D��"o��^M[��W
�\G�����XM&֫�f�8Ɵ�����{�'�Ģk����uwdV�n�
aI��񬊒P�7OJ�uyj0RV���S5�BzG��ӝ�eU��X��/�i����LL
�`p'u�L�`��ەZ/��ͯզD�;t�����/��`�j�� ��1��dk�h~���B���§�I�2r�?�d#z�R�Z��z���By�I^�b�P��p)� -p)2/N������ ���D�9��������Dn����I�{7��
'h���F���+�`E�vO��rU�Ϝ6��nJ�3Ɣ\7����[k�/�f*�l(��3�̱�&��ASTa8	����v�5J��/�Zqڡ�A3B�'������D���G�x[r?�9Z��qU��x��Yߤ��ϦY\��٩ �E���z���3E�[K����\w�q�;.�R��6�/�{1��z8��V��ϰ��Ǻ3j�v�9v	x�\p{�,r)f5i�3�D���Tm;Jk_
0�w黙 �#�5����]>�U�R��Ӧw��S��������8V����*�T�g��3��<���L��}�rŤU�<<�	mK+7�r����:5�2��sN\�t�(�1HF!K��P�y�L�zٸ�(\�b���������tzf�̌���tG�u?\p����jo����� ���LC�i���
���$�)M&m}v<�X������F�Ѷ{�V�eJi���<�/Q�[F� �PA�����jH��P�N��(�̐����3�Oj����D"��w�|�/�*�2���N`���"� x�ѬXH����=�j��� i��Z�\���gS]&G�Y_���쒀��V���R����ٳ�u�{'T�]y��)����g ��q?<�?�d���zPgQ!���~:�y(8u������\�i����aw@��:q/�y]Z���q�<� ����;�=ֳ@�N G��淀�k38��z���6"�0�9�͆�t�:l�6mu;�L��t�`凉�%���Y��:�u�H�5����0�%�T+�Q��6JN�S�p�YIy�X�� �gm�C*��Q�
]���u��� ��n�de�&�]?�"�Ub��]V/����4u��d�����Xה�.�1�7q[D��v�4�����Wn�)����w�� A:���B�~���S2���Eŭ��/d�0Vx+=�e���?�;WP��8��/TU�i��(��|��U~��>Svd�y�����(�B���U� na�0�1�~�N��/�|���D&���C���kV0��̠O4uUG0����767�n��eKe
��6s�۸�遲� g���coD1l��u���m�gVg���b�:^�8¾�7p+D"'gG�/��I��K�Q�S�+;u�T/�r�$�X��A��|�񧿬p� �U�^�k;��� *r�5��ߓ�*�s��ǽM1��y��9PHg�3{�4�����^c"�1T.��#V&�NJ2��H�:���y��ըE��~��+�P��Q�2�C��zk�E���������͌4��nο�p �Vv��i�C��~�Z(��[9�}�z�o�K+��]әip��{��2�!�_���A��jr�%Ȣe:h4F��J�u��>�q�$��1�KG��Z�Q��0�*�2��b��"�����O�\���I�kML���O�I�.�!E)��+�N�������q/��*#-�=F��.	aH=��#!牭y��S�bɦ�h���J�"x�0H�W}�1�m-ɄrIK{o�eB�7{�O�?���&���J�-?236�D*��kC��jm��D��Bcpa')d2<:�j(g9�B}5�15�Ϫ%>�A�<P�@]�8��-!���.I$Ǿ�^�1M(�������S�J��q]�w�H~�[�T��8���=h?.�"�����E���l�맸Ȝ�0��E�����0�M'��ȵ�4:nz�ג�H�m���2_!%���p+�![��V20��ٵv��2���!�8�7��<��yě5�Rw#bz-�w�.Y��\QuT���#��b-��u��IJ�ҍ��AT�2V�����W�	̞�A	�������'�d=˳D�L�ޗ{9��x��qz���??f��_F������TUrDz���t�,(߄E�9q,���å�mM��
�a���ѓ�m�sqT\(XRl�����1���y�DXg�\c-��e�1rK�5^��>+gg���"S�{{)�D05��+��<E��d���|�3-�9���ݽ6ª'�ɫ�j�������GA��f��fB�����	+�-���=�_�j$�s�<ڑ�7p�}�	 v�ϥGq���3P�5�q�0�����8�ـ�����
m�J3Ig�= K�?yJ�Ʀq{7�������ru��cP�� �����M~jW���=��]���
{T�4�$�9
�Ff(�l�]]����1�`��c�y�fd0j�c��P�'瓂��F=/O�O�S��*�
+㮘������Y�JG���P�j)A�J�S�p��q�a�tP~&��v/���Ĥ*��r�QS3,F�8��ĭt^���]��}��N��0�I<,$Z|ښ�m (9�cx���uK� ګ1x��j>�"�M�%��mR�ށm��]V��aҶ��#�K?Q�����թ%Ǜ����R٤�Q��Q�#���ꍹCk�(���A�=/�Z�I�z�<&��U�� �WM�>����e��r��R��]$�Վ'̷^�o%������ ����=3���
ߏ
���z�-���d�����B���	a����@�;�ʥ\O��Ű �M�7��,�2�(Oo���z��7��$��@V�Sr���Y+=�͐l�`��v���K�U\;�q=-��P��=�����S��h�Y\��	�c
Af�Kd@�����̳���ű��;����Z��܅�m#���Y\ȟ�J�ѐPlS��	*���$-���)T�p���'K>��
<RKD.�"����V��h/oB����x&+���i���r���ڌ��Ỉ~�'�R��8����4<�k�5��޵��4�N�x�	$�D��g%���Ԗ ՗�Jb��
S�iuɽ4*#y�)i��֯���t���j��g��؜8�� Z��I�qL�V�^��Wq��9�3��:��21�I,p��7djp�?]��U�������;��q�gR-�A���|=�/�ɃkE[%��Ʈ����m������&��T�05l}�ۘd�g��^����u��0�]���2[3��u��{��:��A9�r���}ު��X�:�>iL��.Y�;��v���rB����n�p��&�T��V��W�����2��������X�<��D{m�.���-����B4��8h��V$(mia��z���x:���}>r����_�\ЌR|ښ���M����;��lKXghĮ�*�gi���X_�9�ߟ�)i��!����L�h0��W����g�?]:�|�|��!�EDFJE��� S
y�=T�܋�����l��H��X��t��YG��`j)��r+�Lm�.u�Ü�|�;(�E�=�Ossg���>ul� ��������������0� M̽rNּ���Lc$-S7�����2p,R���P�N��c�S9��5B��;Pݸ�k������t�h5 9m76��?��D�}���^H�B�
���#��j?}�0Mٿ��� $�SzP�C�;H����X��X.�<so�w�������ʦ��O{w�����7��e���m���͔v.��њ�)�!�� �-X�B���j�Ѓj����,����Q,�W8$r"��а��+DA�/?&~�l)�c0�%�It	8��~e��m�|+)a������uyIS���@�֮�G"�C@-A ���\u����eWb��@���#B �Z��y^�,��ц�>��ڶ�ܖ�?�A��H[vsȷ���ʑ��p�ĥo��㰧�s�Jm��2�D!����4�j�a&w-�̚�P��9���p��N�&��<`א�F��?���_��s�Lc1���UޠEF�s���w���*=chcPt,�L&�0{�"��X�CcU,ZPIm�j`:B�B�اQ<������������١a��5��&�r�@��@�X�	��o�����	9��G�Yc"�}������97�-K��4ٚy�R��wCi������J�����0̮1�j׌œ���@G(�{ZAR=R��ia6��ͻ���"S����t"�=��Зe /-�>��!���en�D��3��]����lq�KҘ�7�]ٞd`�7�~< ��7��rnrw@���)#%��O��+��KS�#�[5��K���+�B��xI��5� ̉�J'�s�0�D�Φ	�s#7��򐐘����k<dR �e!���(P~���?՜r�d��L_���w��D�d�v���Zs:{<� 䞍x���h�l�j(y��o_�l�4w��M2�]�3�3����I��K՜�[�H��-���'b�j���h����暳j�L�\?!��ܒr',ѹ�$p���8:\_K���-ӊ��a*:"Q"�7�a�����"�Y.M ��L�U)�O#>!�é�����0���J� ύ�?��|�jIv�.�@�å� ��!sT���WR�W�<�c�{
[8|�A��k+jm�?x�ձݕ�̺�M�����]�Er��! �?����p���OBW��ƳĚ� u3�?'�B)T#
u�~�x���R�m���}�J�I@�%�o֜��1��(�%-7-�0ůe���$��/b岕�	�s�N�ۙ�����Y��*R�:D_jEJ��_������8����e��p�i�2C�L�K+˼��H-���GqC�F5)� �=ɢ����_���D�jJJ�4��Ԁe��<���ܧ��$�Eu^z��YǠK�$'���Y��t(���U*�1��`?B-�H��1y׿�7�+��=���sp�-�Y@C������D�<)�9&TaN؆�l�X�0<֮��wN�_M�D�WEV�����u�܆�D}T�`}��Ѵ�S�����c�e�\�q�q�������L�T�S��!�yZ�n[N��������sE]�D���#��b@�3 ���~e�`l+δ�A���f�12���k��<-@_:��[���_pa�m����f�h⟄ᨙ�G�~R`%�Ő��>ָ��(��d�>Z?WK�IJ<m��b�鷏퉗���L��9Sܺ.K����%C�5��=�ܘ^��|B��)[B�!�*2T�%�TS ��.Sx�:�9��A�g�]v�Em76��;� y�U��p�q1�V�6���O��7{Fh;�.3����@�Q�s>u0�vގ��x;,��U�]�u;jUP�X�B�n�)I�"n1s��ZK�!������p�t�C��
���^V�[�d��U;����N#^Y�ѾGS�!�)��G�d�M�3���/k<c,�r����ښ/�hٹ6�p;&������}c�|u(������OsXC�6f�M���#\�b�:�U�>~����9/�����$�َ�7��\4;'�ct[�DVl����	�o?�5��)�8l7>�$W&��k��������⎀�=��M�NG����0쁇�'�e�1G��WϷv`�H�&A�m�W���+;��&i�fA�T�os`���$�,��j�.{��!� ���+[�f��pyy�̘���wJ�9TF�"p&�������Ҩ��j� �7�߀�	Wq���c��"�Ŝ�/����V�q��e�|��s��A��Zи>���5���T��;,�Y���>-��D�XZE�����X���ׁ��I'���P7y'|\�|�@�ԪсB�l����﬿j"s��T���c�<��^p�){�!|�jP���1S�V���'�ؾ^p3xOmBj��mP�U1�%͏�6�_�^O��c��.k�iC��љߗkq|�ugM9lJ�����¿.�'��Є@�R�j>�4���m���>
^� �����]���W�*,8�v8۸��*�V1nFz�*�n�>y=������	��G�&.�XP�W�p�b��7��i��Ӽ}��Nh3T!q����=�ui��:��Gk�e����v}�Ue�A���r���@#p�(|���p��t����$�Ԫ-�'.?�in�U�\�{H6G����G+_K )���X#�)�x].�o��X��ٶ{Y�Ѓcq �*f�^qj��M,�ׇ�B,/��󼩘#�p:p)l߱�koᓉ�я�c)�+����Ɠ<b����y�n�����TL���%#:W�Om�VPN?2t&e�Pmŗ�����)J�|�#�1��9�Z8��·��#���y
���)o ��©a����߻�.�JO[��77��Ŏ���+|�Җ�"������6 .>�� *
k�(�Z�[>/��/�7�L@j&�q�T�Ua�/�`���|s�,Xf�ҿmƅ���A��X����@�8�fb=��a+���tp��Ă`�|H�S|/Ql4�\L���Hö9O�y:O`�{�ִn��;ȳ�T� $�Y�E�S�Wg`��f��-�=��r��V���h�6�s�2��աSr�1����y�X���^$���/pqD�I�=Dj?��|�!OA�*�n#���L����}����'�E��ܑ�����a��b�$S��T=N̈D���S>�1��� *%a^=��U��g�>m�5�w�tE>
�TO)]�i�*�%�}Ș��u�-5�8�S6�y���Sl�� ��ۖ3hu�\����H"���"�X��*-���"�$��z����_-�轌�o�I3}������QiY7�x>�l�_ŀ���u&$�d�D����f�X���CDpΞ�C�T\����9�|�ڞ�wTc]7,`���a�J5t4կm���a����T��	Ut2���D�i��'���M�� �em���`?�#�]�b���l�3�L )���(3�jG/%���Ѻ�j�́6&Or��ǣ*I�& �ݮ}NΝ�>2_�_�}�:�sk�y��=3og|����aأtokum��E,Ad����/6$9e	hј� iq]	�'�^��h�D`ŝ԰�9[a�bk�im�{�7��y�#���I�u)����g�Y����Ǡj_���keOh�Q��@ s^ƾ��1ʬ�&�����E��4��p��ƛf\�،l�U�l�*���$����6ˬ)ݰ�L���M�H�Nz�t�TR����'4�Q����l$wNZ�$�7Ǝ���@�A��	��2�:�:��g�i�R!�"����џ��H�g��{���:�3M�B��T��,�pd��,4�I5�M��q_�ֆ���)�t��K ؄`�<=�ݪ9�� ��0�0�I?� �%�U���4S�F}�[sg���̌�"q�h�JA_߱C*��)a.�ΐYK�U;�G���r�q�c�Ș�oQ���T
�����᩠=8�!��e� �u?.�:+3nV�E*����|�b�W������|���QLv�2QH�PG�����+��&�ລ��;\�Q(��L�a�<]�I�0�*m��7�z}ċ��8x�	i�k
����TG��>3� �f�5f����/C�g���L�� ��us�\�-FNO�s��ŵJ4Y����P�m�ds����Jr}1�R��$�h:%����/��-��
?���

����KX�`4�X��o��)�}���)m�f�^�c�F�`Ǆ���o/鰯I���pq�1��꩷Sk2$�� ��,�%�����&��3�)�@�E��x�c~(7썋��t���T��=c-B��E��S����Y��P���Py;��[�,�l6�q�ሲԮ|^t��Z�.X�&��tB��>�i�� >D�@��>Dv��e��V�pʬ-�/�����x��ы.Wj�(Ϊw�a���0��VcY�.X\6���5y�j��3���}A��LJ�-Eڠn��~_E����q��N�gߐy�X�,s~\�&-����xK�p��7�Nރ�ր�	��ڏ��j�x�8T-��јS���&�Dkm2�Aq 1Æ�W?�S�����Ӽ�9?v���f�����{����~P��qw�Cz�G=Ԍ`���C@�����OBJ`�� ���#��z�o��f�eH��Dk%G+�7����c."�31F p�����g�RP���'���7�DG�s�Oq�o�2� l���;���@�xhJ� N�pjG��W�F'���T?C��.�>��N��H�}�[�j_Gk���SH�v�!��5i\Cs�F��i�ݷX)&�ob���tfe�R�$�`��G\�a�.AF��o�h�t}X�^^���]P&�q��h�Ke*��fJ�cn���n2@7����]��8�:F�ˢ����D��|� �W!�x�ݎ�x��rٛ�4ex��(,P~R��8���w�"������)�#~��)눢Q� �t9�W�[6��|�hZ�A�N�
˅�*3��y�D�}����׎}��)�< �I�Q��%u����T:�������䈇����p�٣p�ٝv�p�4�&��(�I*=	mn�W��̲/�wtQ��e(Q3��l�~BS���g�Wd��������3�4�^�;-)�KN��#!W�c9Rt��rʬ��2c8*q.|�kf?G�p�.Y98�Uġ�` 5�0I��!S�(�|�����u)���W�*����8�"T�#��*�Z:�S���qs+ T��&��F����g7x�>?N�rG��|S��׾[�(��M���+m5��V&X��t���9^:#�r\;�˾�u(q񅂦��f[1�K��K�B?O���F/���#�4��������|uIG��׼�|���C߱s8.��p�id���p��=-�3�P�4%H?��
���4���C���kg��s�C���[JDu=�g�~,`j�|Z.eH
_�٦�j�7�o��g�i�]�arnB�'7O�Ȃ�ׁ/���1���]j�|Q�_�S �T�"�B�S�ޜ1)W��SΑmGg_�����3!�����8�2���5�N��s�'��"��hn3��u}x	�q/X5�b6W�и�&�1˼�]����A��J�Z:�>z�XE��I�BU�_H6����A�;)Z�..�5�׏"xr�����>�kJ{ϙ��e��)Es�d�]�n�oc��⎵��$N��D=���j�zΘ�{��n���|�V����A�|` �k�;���!#�l>��M���S��3�]!$X��@:͆!�u��Ա.���&>=����ݩ�b�5�W���E�Ĵ�x۳R����\e:�C�����ň���`Q� v��OCƣ�h�M�f�b!��(��״wO�XR����^�[1o�#��G^L�x��`���ÊN !�XD.��0�@�li�GM�������m%�'h�m;+0� YAG��ԟc�<����H�����K�7�����j�����8"�\��f��78?���X�I��*�,$%[d�a�^k	~[����h�a���Qq���RNͫRu2%vY;��*w�9��Wh9X�0f�U�]��͏3G	�KrDie�+��_�b� G,��a�n��/{�CHOI�߫d 5�*�l*�&�����D(�N�<5}�ư����LSxr'Q���[��u�k���$ꕆ�&�u�cSZǡ��74w�J�Sp��/��Ŏ
C}�BR��@�A���9��٧.O�S�1��2��n�"���Fwr�{��ߐW+s��p��3�L�
��Ȯ�����i����{ӌ��A�r���wF��1�x^�!K���*J��8�V�xbl��i�^] R��MB%��*@�d���C�/L���0PFL��JHv9��f����YZ���]��ν@;GS-÷�=k�Sb>Ȫ��i���f2�}Z�F�������s��թ���s+���hU��Y&�c�8��c��OW����ԥm�p$G$� ϢX�\b"�4�'����³���10��ͥs�ӴP�}`�?��';=�gtB��4/�F���^��u �=��@0$X��E�Mw\D�}v� h�hr&1��+�s���<�i<GC�>��"�����H���!�zY<�j��uo�k�ٍ�F��a��,ܠ4}� ��]q���g%ݤIZ�r���|������_,X����3�R�H1̈́�������sy��/��U=�oZؘ��\��t�)�^���m!���m�,f�ի�A�Z$����٫?˫Y�;���G(V�	Zh�E���o�Z�y'�w*K�@�a�.��r�Eg��si*�u?�D�F��-^�	�4��Cd.<�gW�k���v��{��8�|�kq6K�hgG�A ���h�E�e��{BBO��F�����e��'�+�k��y�
�ީ�
���W憊�Fł�%[�z������m]�c�:/A�S�e4��.qx"��N:2���9G��d��o6�l3pV���~�V��.jp.zcy�$S��DP��^!ʟD���f1��;��|ly�N�φ�2@�*W�lafM�L꘲V_�*��4�s�ɴ8��o��D`���y�ϙH��+v�T/��7N�ɼl��%®4�60j��j��(�%�!|���lB;iňpN����5�_H�5#>�V��W���JH��<|�����/u��)pGܨ�+פ|=m�0�.j����`;����	6D�Bui2>���E�X���m"r����qZҲ䳹k��^<V($��;Y�.���LL�Ϫ�fx0��	v�vXN5��O��/)�ҭ9Q;�h������QM�t����s
0��q.�3����2�$�����C��<�ʔ�~P����Xw�.51J�tH$�w`Æ@`;���`b<�޵�X�Nq"Ŷ���[�� ȯ�EB;ϳ&߳���u}�L����+3$�Ӂ
�oZ��bX+e�KFxH˅�f��]"��'kZ\�ӗH�]����Y;x���2��ޘ�g @H̾�P%���2[�tÆ0��C]�!f;z��V����"�t*ku����~�sz�zܣ�%�_��R�z��$��o�{���ٗ�8\I��:4 ��/���4���'�k��*�g�y�̳��J�Š�7���M,�ae�`!Mp���r;�i��~dk�>k�	��b|��{�0�Eՠ�XNDЍ9}D��y�Z�����(�2�)L�>���D�w�����t P|6���Gס�}h��3,���ԫ5������/uMB1=H"4{����}Y��,�Qb?��kw�E�e����[tMS<.,��[]+ )�Ӟq"�M;�.�q��+�φ�Y��+�OA�`njp�}���(���~� ��TĂi��"��%�U�_��S��7Wc	�:KX5������	���2����CxQ5>|fє
������R�5��ї���}kK �* e�l����cS~?
z�z"�[Tj����ژ<�zR�1���q���OQg�~�(d�����3|ٿX�ޗ����2,�8��$I��~��|4o��$�@?���k\R��3�3�YJY2귶�������v5	aeD�#{ *�����f"=:G�9��nId�K�fVC�ځ�kMU����YA�U����_�U1��8�qB]ԃ���Z��ȳu�j��,��?Z�1�;N�)d/�e/��XӁi*��+��"��4�8�`�� u'>D����Vmb#��Vͅإ���6+��#��zEq���O&�؄ha��=��q�+T���(Ȥ��P����f��6`��]l�?�=�岶���u��T暶�
-j<�4���2+1
a�f���d,�q�Y[�4�q��gj��{�B��'�-ɟ��Y�6��D�h��P�{�l9;b��AE��ؚ4T�=�-�2؉����a�0oS�5� ��^~;�y%d8:m#�V�/�c�05��H�6˾��Թ�k몸;��7v]<ԩli��[EZ��g�f,@�Jf�>]�U�����Z�D��[O�87=��9�3U�#ga4��Y���^G|���_����C1�Q^�w�3��1a� GL���uR'�ok>���x�\��هH����}zz�=���!������Is��E�����#�|�:�-#��?���ή��J8������i,F����0�RX�;�=M��^�N�?l� �_�A�j:�1Ѫ|�}cp�[Ǆ4�.�0;����m3�/!��B��O	!);[�!� O�����XmB�<��	�c