��/  ���T79'@yV2��:T!zf�g͟��a��WI�s���%퟊�e�c�\����[�t����j�X�8�����$4L�������}g7l�� *��I������,0�z8O� ��t'�O��!y}_���C���cC&��BB�m����_�2rI~�K0�HR3=�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC. �,"��'��g�	���:)J�U��>F���\(V��S�Y0�$�Sv�ջ'�c�@��mt+�:4�.�Y��X\
��z*WR�||"�i"�����ᓇ!�I+��_�Ph�5�5&ig @���bl����4Lꭱ�jy1Q7�r\X3p �Y|���u	��[e�Ƕ����+Ƴ�K��$[{��ha
����6�{/c�wD��J��R, `�s�K�7W �fr�!o��;b���A�ͺ� ����\��o�XŖ��N+�}j%j��O~m!�׹еv��>�r�6������v�� y,ۆ�]@}�:�e��=���I� �~��czK�PB��H���z8H6��7R_&�2�m�Z�tܷQ�2%��C�Hf '׃O_ځa,�ؤ�<3~.;|J�R	�j!�ld�p��FtCo35a)���vډ��q����J��X�h;o�/� އ>m��J�q4A�Kh �{�Q���4j���<���ǒ��L��V��!�$y=�^�v&�ī��� ����\4U���V�h.�/�,];���&!1^��(N;�gC1nǦ�/�4�e�L��f!�Ao� �ŝ,gq�r���QI�Ū����Gm%�n���ܭ>A�H��P��JLEEQ}�$6R
N�9�ϯ[��c���ZtIe�g���8h�{m� I�`6
^.Ya�V� !�Lе�B���+iu�N�Ρ�x<�ѓǞ��� �%�-fgk.�D�o��*s��}%�ػZ��iq��?0���'�ԭ�$(cF�����+Z�i�R)��T���n���E�����/��F�[�� �4����W໪���j��<=�1S ƥ�ofR��&H�)h>���c���);U�GAtR�R�>�u$��9�|�W�oD��G��9�O[�����;�ޕ�u�U��ߺW���򲢲``��UtE�^���؈���k��
'[|`�a�{I��.KƊ#X����ʳ�Z~��e+I\�8%�E/��h�|�)C�a�p�?n�ˡ��8�֥���Ny��М���x#[9�b�[��=g�C��}��4Z�}*��] {h���'�Z�@��ݜ��@����Z��4�m�ږv��r�s&��y�CZ+׫��<4�������?=|��O��-�#��@����oZ��r�c7Q�d��3u��<�0��+�˃P�I��[18\k�9F[ǫ�J��T p�����,����� �м����(����»�tm�2E�h��^���y��v����3j;ʇ����A�Mp���3��(���i0H8�=�vm$﨨�ё���e)Gs �}�Y��7�m���y� J0a�L�4�+��3r�'����~�(]*n��0>F+��q!��{�i���"���9Re�F�_� {.W"� ����M�$+����6���DӦ�b�zR��H�七�� #��� O�P�A�W����X�i�O�H���m5�����u�f���F;�n�����sC^dX��O�"�^� ڦY��?�/�l���O��H\,aFo2O�NWd}���G�f��G�4u��)������
B��D�r��]�m�bV4���uwE��@��V(f�9`���Ǿ$�΅��|K�]T�pna��.���|��Y�t�A	��z?����zg�5m=�*殇����oh�X]h1+��uo�$����a}���0/㘬Q�{C�%ڀ���D�S-�)��.Ĝ�V�B��)\PGp2���W��H���"��1胤苃��E�w��A����;���A�v��!׼E���d�߁����8�N�p����q���n/�n}����aě=���}�z�K2B+�⮭�~��S�F�o���}/�6�2PG[���r�/}�?�	u|��N�O|��.=���zh���\��A����\v���/>,$A:̿_"�N�����H�*2��k��le8ӺM�dL�l��S��%R��>å���7��t�<��m�|3{w�mFvb� �$��9?�5Yv�1Vg�/u�笨��ؑ�V�%�a��|W��9��=�)á~��0��V�Ko`M��������+�zvd�Q��M�!�;�jr�\�Ǣ�����BwR
�Z����}�����A"=���HE7 *��-�Kd>2)�!E����k������	���0	�v�k�!0��	�{���������0p>�ټ��?��⯻ɋ�d6@U�k�	�9/h��ՙ1�,�gp��/����6�\�ώ��o��p���7_����+��,0��N'�DD�'2 /�D\�|���1x{-�PI��ٗu����)��P��jW'v��B��u��.g��r�!��LS�`C��ͳR�F���M��b��bb��h5�l� ���\�0<Wa;�P��F$�>��_t���)ë�)9��Y��D^��j=�/���U�s�R��'S���S�Jn�(0Yc�����1�?�fPl���X���i�Wc|vGP�[+d<�ЀkQ�=�-4u���è��+ی��R�la��x�� ����L��ʀ�1���Pl%X�����Y���( ؖ�Ӫ�]x��{@(�fi͖���'�ϒ�����ֿ�T�9�?M+��7��dt�؂��2@QQ����ϛOg�t���iJ��뛫-�˧tz(m���_]�+��~�eD��h֣R(�I����p��B�Ks�����������s��(�<՟ɓ�8K<���*�Za������0�t�qt�Σґ����(R1��JlC�d�泌\n�%	��"�9� �Lb�*e.��.g"��i���@�p|���v�X&�,BD��R��ƜE�IVA�-OP�x���a�nOw	�]r<�ڪ�������K���	
�I�S��Q���/���#�L@ڎ���C��k.j�{��%�&^Aҥ�����P�4���A�|�M����j�s]yR,,�c¤�T��ğ���q3�%:�ȖX�H�.�Ԗ�1����J��X��,� )�)����;���ڲ�sh�ݨI�/6�l�W,���)��L�{+(�[��$�]�OGD�q����/ؾrmo�fg����|3�uX�UTYV_��O,^#��J��wo+�����ȯ(Ȍ�ƆA�4����<mh�G['�,���1ȂWṑCC�˾A�xp�-�ƺ�I~5��˗����W#o/J�\mt�]*�2^���V3�?����M��v�>7�� �c-�
�����GtY)R��y�F���2�\Gӂ���{�]	Ul�,�؈7�y�\ȭ�G�V�����1��נ�"�R�~t�[T�|ދq��Q��� ]~���ec�1z:�!��9Ʀ�sS��(�2B�$�A��n�-P� '-.8�۸���_J�|nY�^?�}5}b�a{ dN���0𦙞q�Y˹V0��[*�]s}���?�~S��xE�5_U}rƤ�	[�`"� �4����ҋ�������V���K��e��PvW5%#�G%鮖K}22��ɦNCzt�����`���JE�6��W���*��/4��K���dS_A'��4�)N*&|s�º��w�d���MŐsl�u�)Z|� �����a �?������K�#7	N����Y:Q��1�	ݰ�*�΍�s7��x������ AwO˭��|϶ڧ�\R2u�[�<��	�P�r���z[�sTiS����"�����H�F�~5�9#���/�v�'��*��n\x^#�#����\�i�m{G�`j�I'3�g\�4Xy�Z���)S�{��B!�@�-?����y��O^�Y�Bu�M"�x���G1�<RN'~��c�����B3�7����7f�t{��!�n��VA.¾�.p*��><���bJ�U�Х$!^���dk��VH�%ѻ��B��?��?A,?��z��˄�c��,mc�nK:K�}��5��f\X�y�j͉y��30�m��G�f���=h5�58��/�v
�uuG�l�9����ao�/X
�*��Jl�)��HL�I<���J3Y������q3�7-Tכ�k�!�_�����I}	���aMi9�uW 4�[z��;D�"&i��BL?�z�N��i��ۀF:�Z�@�x�!��[g�.~ �B�9f�΁%B�������#O��:t���s�%��lUÝ\:%:�m{�"��W+�]6�Cc|���<c`'�=>4�W
�����b*�7�6+��	��+7�QojmQ��U�q�I6_k�����NR���V��1�Pά|�ù݃���2��DZ�j�ѕK��*�8_	ރ�{�����@���B���ٽ�g��MEl�2-f*���ھ)p�~����ئ!����^��'��+Z9�ʈ=^u)��}��E���o��� m��zv�mn��ꑊ��h|j���^U����/��m�X����78��6*o�-^��p�@R:���T_��� �Gr�Ǿ4����(	��,ěeR��i;����M@�"���
�P��έQ�Q�=�YG
�������54�O&
"���[�γa�=���C�U��A�	��c��=%ln�XB*���
�q�ܮ� P߽��W�~���!�Pn� I2<�
֞�@O�F*t�s�|yT�!e��[�!~?e\/��y�HD{��,G����b�U+��{�NcE�XK����j}��sO�[���{V���k�����JC���a3`BO��&4(��Zw��ˡ=��p(?�1����MΟ
�*������%3}�*��.VU_s\,q�`�>�����^��Q����x+9���b}e�wخ»	\-���e��D�؅����jV�J����]pK5-q�_��tyч�}�3]E� "GT�����y~����^VUu��n�TLE��+Q+�vI�a!\Xw�\??�-���]Ų�� 	$^��"I\�,D�����]X ��ek8�p�1V�O�+ �%������S� �R� /0�&�x�T0q�Ra俵D��_���̵��{��I/�������@Ir)V��9
g�9'��!�	ݣ �DN����E.'��V��fl#��/O�t>��ʬe
��p�R)�Fh�-�|:x	}�z������|�C�q����4P�a�^Y \��?���pb�'�<. �2��>�����d��x�9�l8�wo�7M���$��(��K�S�K��V�#�o